
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE WORK.pix_cache_pak.ALL;
USE WORK.pix_tb_pak.ALL;

PACKAGE ex4_data_pak IS
    TYPE cyc IS (   reset,  -- reset = '1'
                    start,  -- draw = '1', xin,yin are driven from xin,yin
                    done,   -- done output = 1
                    drawing -- reset,start,done = '0', xin, yin are undefined
                );

    TYPE data_t_rec IS
    RECORD
        rst,wen_all,pw: INTEGER;
        pixop:  pixop_tb_t;
        pixnum: INTEGER;
        is_same: INTEGER;
        store: pixop_tb_vec(0 TO 15);
    END RECORD;

    TYPE data_t IS ARRAY (natural RANGE <>) OF data_t_rec;

    CONSTANT data: data_t :=(
--                 INPUTS              ||           OUTPUTS
--  rst    wen_all  pw   pixop pixnum      is_same   store

	(1,     0,     0,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     11,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     11,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     11,     0, "*:::::::::::::::"),
	(0,     0,     1,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     10,     0, ":::::B::::::::::"),
	(0,     0,     0,     ':',     14,     0, ":::::B::::B:::::"),
	(0,     0,     0,     'W',     9,     0, ":::::B::::B:::::"),
	(0,     0,     0,     '*',     1,     0, ":::::B::::B:::::"),
	(0,     0,     1,     'W',     11,     0, ":::::B::::B:::::"),
	(0,     0,     1,     'W',     3,     0, ":::::B::::BW::::"),
	(0,     0,     0,     '*',     8,     0, ":::W:B::::BW::::"),
	(0,     0,     1,     'B',     4,     0, ":::W:B::::BW::::"),
	(0,     0,     0,     'W',     5,     0, ":::WBB::::BW::::"),
	(0,     0,     1,     '*',     14,     0, ":::WBB::::BW::::"),
	(0,     0,     0,     '*',     5,     0, ":::WBB::::BW::*:"),
	(0,     0,     1,     '*',     4,     0, ":::WBB::::BW::*:"),
	(0,     0,     1,     '*',     14,     0, ":::WWB::::BW::*:"),
	(0,     1,     1,     'B',     1,     0, ":::WWB::::BW::::"),
	(0,     0,     0,     '*',     6,     0, ":B::::::::::::::"),
	(0,     0,     0,     'W',     3,     0, ":B::::::::::::::"),
	(0,     0,     0,     '*',     5,     0, ":B::::::::::::::"),
	(0,     0,     1,     '*',     9,     0, ":B::::::::::::::"),
	(0,     0,     1,     'W',     3,     0, ":B:::::::*::::::"),
	(0,     0,     1,     ':',     14,     0, ":B:W:::::*::::::"),
	(0,     0,     0,     ':',     13,     0, ":B:W:::::*::::::"),
	(0,     0,     0,     'B',     11,     0, ":B:W:::::*::::::"),
	(0,     0,     0,     '*',     0,     0, ":B:W:::::*::::::"),
	(0,     1,     1,     ':',     13,     0, ":B:W:::::*::::::"),
	(0,     0,     1,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     14,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     10,     0, ":W::::::::::::::"),
	(0,     0,     0,     ':',     7,     0, ":W::::::::::::::"),
	(0,     0,     1,     ':',     7,     0, ":W::::::::::::::"),
	(0,     0,     1,     'W',     14,     0, ":W::::::::::::::"),
	(0,     0,     1,     '*',     3,     0, ":W::::::::::::W:"),
	(0,     0,     1,     'B',     2,     0, ":W:*::::::::::W:"),
	(0,     0,     1,     'B',     9,     0, ":WB*::::::::::W:"),
	(0,     0,     1,     '*',     8,     0, ":WB*:::::B::::W:"),
	(0,     0,     0,     'W',     9,     0, ":WB*::::*B::::W:"),
	(0,     0,     1,     'B',     10,     0, ":WB*::::*B::::W:"),
	(0,     0,     1,     ':',     6,     0, ":WB*::::*BB:::W:"),
	(0,     0,     1,     'W',     2,     0, ":WB*::::*BB:::W:"),
	(0,     0,     1,     'W',     0,     0, ":WW*::::*BB:::W:"),
	(0,     1,     0,     ':',     11,     0, "WWW*::::*BB:::W:"),
	(0,     0,     1,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     1,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     9,     0, ":*::::::::::::::"),
	(0,     0,     1,     'W',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     1,     0, ":::::::::::W::::"),
	(0,     0,     1,     ':',     6,     0, ":::::::::::W::::"),
	(0,     0,     1,     '*',     4,     0, ":::::::::::W::::"),
	(0,     0,     0,     'B',     14,     0, "::::*::::::W::::"),
	(0,     0,     1,     'B',     4,     0, "::::*::::::W::::"),
	(0,     0,     0,     ':',     12,     0, "::::B::::::W::::"),
	(0,     0,     0,     'B',     1,     0, "::::B::::::W::::"),
	(0,     0,     1,     'B',     10,     0, "::::B::::::W::::"),
	(0,     0,     1,     'B',     11,     0, "::::B:::::BW::::"),
	(0,     0,     1,     'W',     6,     0, "::::B:::::BB::::"),
	(0,     0,     0,     'W',     4,     0, "::::B:W:::BB::::"),
	(0,     0,     0,     '*',     2,     0, "::::B:W:::BB::::"),
	(0,     0,     1,     'W',     14,     0, "::::B:W:::BB::::"),
	(0,     0,     1,     '*',     7,     0, "::::B:W:::BB::W:"),
	(0,     0,     0,     'B',     3,     0, "::::B:W*::BB::W:"),
	(0,     0,     1,     'W',     6,     0, "::::B:W*::BB::W:"),
	(0,     0,     0,     'W',     12,     0, "::::B:W*::BB::W:"),
	(0,     0,     1,     'W',     4,     0, "::::B:W*::BB::W:"),
	(0,     1,     1,     'W',     6,     0, "::::W:W*::BB::W:"),
	(0,     0,     1,     ':',     4,     0, "::::::W:::::::::"),
	(0,     0,     0,     'B',     5,     0, "::::::W:::::::::"),
	(0,     0,     0,     '*',     12,     0, "::::::W:::::::::"),
	(0,     0,     1,     ':',     5,     0, "::::::W:::::::::"),
	(0,     0,     1,     'W',     1,     0, "::::::W:::::::::"),
	(0,     0,     1,     'B',     8,     0, ":W::::W:::::::::"),
	(0,     0,     0,     ':',     9,     0, ":W::::W:B:::::::"),
	(0,     0,     1,     ':',     0,     0, ":W::::W:B:::::::"),
	(0,     0,     0,     'W',     12,     0, ":W::::W:B:::::::"),
	(0,     0,     1,     'B',     0,     0, ":W::::W:B:::::::"),
	(0,     0,     1,     '*',     2,     0, "BW::::W:B:::::::"),
	(0,     0,     1,     ':',     15,     0, "BW*:::W:B:::::::"),
	(0,     0,     1,     'B',     3,     0, "BW*:::W:B:::::::"),
	(0,     0,     0,     'B',     11,     0, "BW*B::W:B:::::::"),
	(0,     0,     1,     '*',     15,     0, "BW*B::W:B:::::::"),
	(0,     0,     1,     ':',     3,     0, "BW*B::W:B::::::*"),
	(0,     0,     1,     '*',     15,     0, "BW*B::W:B::::::*"),
	(0,     0,     1,     'W',     7,     0, "BW*B::W:B:::::::"),
	(0,     0,     0,     'W',     2,     0, "BW*B::WWB:::::::"),
	(0,     0,     1,     ':',     13,     0, "BW*B::WWB:::::::"),
	(0,     1,     1,     '*',     7,     0, "BW*B::WWB:::::::"),
	(0,     0,     1,     'W',     2,     0, ":::::::*::::::::"),
	(0,     0,     1,     'W',     4,     0, "::W::::*::::::::"),
	(0,     0,     1,     'B',     6,     0, "::W:W::*::::::::"),
	(0,     0,     0,     'W',     10,     0, "::W:W:B*::::::::"),
	(0,     0,     0,     'W',     1,     0, "::W:W:B*::::::::"),
	(0,     1,     1,     'W',     1,     0, "::W:W:B*::::::::"),
	(0,     0,     1,     'B',     11,     0, ":W::::::::::::::"),
	(0,     0,     1,     '*',     12,     0, ":W:::::::::B::::"),
	(0,     1,     0,     'B',     11,     0, ":W:::::::::B*:::"),
	(0,     0,     1,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     1,     0, ":::::::::*::::::"),
	(0,     0,     0,     'W',     15,     0, ":::::::::*::::::"),
	(0,     1,     0,     'B',     11,     0, ":::::::::*::::::"),
	(0,     0,     1,     'W',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     15,     0, ":::W::::::::::::"),
	(0,     0,     1,     '*',     13,     0, ":::W::::::::::::"),
	(0,     1,     0,     'B',     15,     0, ":::W:::::::::*::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     13,     0, "::::::::B:::::::"),
	(0,     0,     1,     ':',     15,     0, "::::::::B:::::::"),
	(0,     0,     0,     'W',     9,     0, "::::::::B:::::::"),
	(0,     0,     0,     ':',     14,     0, "::::::::B:::::::"),
	(0,     1,     1,     'B',     2,     0, "::::::::B:::::::"),
	(0,     0,     0,     ':',     13,     0, "::B:::::::::::::"),
	(0,     0,     0,     '*',     15,     0, "::B:::::::::::::"),
	(0,     0,     0,     '*',     9,     0, "::B:::::::::::::"),
	(0,     0,     0,     'B',     8,     0, "::B:::::::::::::"),
	(0,     0,     0,     ':',     5,     0, "::B:::::::::::::"),
	(0,     0,     0,     'W',     13,     0, "::B:::::::::::::"),
	(0,     0,     0,     '*',     13,     0, "::B:::::::::::::"),
	(0,     0,     0,     'W',     2,     0, "::B:::::::::::::"),
	(0,     0,     0,     'W',     3,     0, "::B:::::::::::::"),
	(0,     0,     0,     '*',     7,     0, "::B:::::::::::::"),
	(0,     0,     1,     '*',     7,     0, "::B:::::::::::::"),
	(0,     0,     0,     'W',     4,     0, "::B::::*::::::::"),
	(0,     0,     1,     'W',     3,     0, "::B::::*::::::::"),
	(0,     0,     1,     'W',     5,     0, "::BW:::*::::::::"),
	(0,     0,     1,     'B',     2,     0, "::BW:W:*::::::::"),
	(0,     0,     1,     ':',     10,     0, "::BW:W:*::::::::"),
	(0,     0,     0,     '*',     7,     0, "::BW:W:*::::::::"),
	(0,     0,     1,     'W',     8,     0, "::BW:W:*::::::::"),
	(0,     1,     0,     ':',     9,     0, "::BW:W:*W:::::::"),
	(0,     0,     0,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     0, "::::::::::*:::::"),
	(0,     1,     0,     'B',     7,     0, "::::::::::*:::::"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     10,     0, "*:::::::::::::::"),
	(0,     0,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     9,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     14,     0, ":::::::::W::::::"),
	(0,     0,     1,     'B',     9,     0, "::::::::::::::W:"),
	(0,     0,     1,     'B',     2,     0, ":::::::::B::::W:"),
	(0,     0,     0,     ':',     6,     0, "::B::::::B::::W:"),
	(0,     1,     1,     ':',     8,     0, "::B::::::B::::W:"),
	(0,     0,     0,     'W',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     3,     0, "::::::*:::::::::"),
	(0,     0,     0,     '*',     13,     0, ":::B::*:::::::::"),
	(0,     0,     1,     ':',     11,     0, ":::B::*:::::::::"),
	(0,     0,     1,     'W',     10,     0, ":::B::*:::::::::"),
	(0,     0,     1,     ':',     10,     0, ":::B::*:::W:::::"),
	(0,     0,     0,     'B',     8,     0, ":::B::*:::W:::::"),
	(0,     0,     1,     'B',     3,     0, ":::B::*:::W:::::"),
	(0,     0,     0,     ':',     9,     0, ":::B::*:::W:::::"),
	(0,     0,     0,     'B',     0,     0, ":::B::*:::W:::::"),
	(0,     0,     0,     '*',     14,     0, ":::B::*:::W:::::"),
	(0,     1,     0,     'W',     15,     0, ":::B::*:::W:::::"),
	(0,     0,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     5,     0, ":::::W::::::::::"),
	(0,     0,     0,     ':',     1,     0, ":::::W::::::::::"),
	(0,     0,     0,     'B',     10,     0, ":::::W::::::::::"),
	(0,     0,     1,     ':',     8,     0, ":::::W::::::::::"),
	(0,     1,     1,     '*',     2,     0, ":::::W::::::::::"),
	(0,     0,     0,     '*',     2,     0, "::*:::::::::::::"),
	(0,     0,     1,     '*',     15,     0, "::*:::::::::::::"),
	(0,     0,     0,     'W',     0,     0, "::*::::::::::::*"),
	(0,     0,     0,     '*',     12,     0, "::*::::::::::::*"),
	(0,     0,     1,     ':',     15,     0, "::*::::::::::::*"),
	(0,     0,     1,     ':',     15,     0, "::*::::::::::::*"),
	(0,     0,     1,     '*',     15,     0, "::*::::::::::::*"),
	(0,     0,     0,     'W',     6,     0, "::*:::::::::::::"),
	(0,     0,     1,     'W',     12,     0, "::*:::::::::::::"),
	(0,     0,     0,     'W',     3,     0, "::*:::::::::W:::"),
	(0,     0,     1,     '*',     2,     0, "::*:::::::::W:::"),
	(0,     0,     0,     'W',     14,     0, "::::::::::::W:::"),
	(0,     0,     0,     '*',     7,     0, "::::::::::::W:::"),
	(0,     1,     0,     '*',     3,     0, "::::::::::::W:::"),
	(0,     0,     0,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     5,     0, "::W:::::::::::::"),
	(0,     0,     1,     '*',     12,     0, "::W:::::::::::::"),
	(0,     0,     1,     ':',     2,     0, "::W:::::::::*:::"),
	(0,     0,     0,     'W',     4,     0, "::W:::::::::*:::"),
	(0,     0,     0,     'W',     2,     0, "::W:::::::::*:::"),
	(0,     0,     1,     ':',     6,     0, "::W:::::::::*:::"),
	(0,     0,     1,     'W',     4,     0, "::W:::::::::*:::"),
	(0,     0,     1,     'W',     8,     0, "::W:W:::::::*:::"),
	(0,     0,     0,     'B',     9,     0, "::W:W:::W:::*:::"),
	(0,     0,     0,     '*',     14,     0, "::W:W:::W:::*:::"),
	(0,     0,     1,     ':',     9,     0, "::W:W:::W:::*:::"),
	(0,     0,     1,     'W',     13,     0, "::W:W:::W:::*:::"),
	(0,     0,     0,     ':',     2,     0, "::W:W:::W:::*W::"),
	(0,     0,     1,     'B',     1,     0, "::W:W:::W:::*W::"),
	(0,     0,     0,     '*',     5,     0, ":BW:W:::W:::*W::"),
	(0,     0,     0,     'W',     11,     0, ":BW:W:::W:::*W::"),
	(0,     1,     1,     ':',     4,     0, ":BW:W:::W:::*W::"),
	(0,     0,     0,     'B',     4,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     2,     1, "::::::::::::::::"),
	(0,     1,     1,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     14,     0, "::::::::::::::*:"),
	(0,     1,     1,     '*',     14,     0, "::::::::::::::W:"),
	(0,     0,     0,     'B',     5,     0, "::::::::::::::*:"),
	(0,     0,     1,     'B',     3,     0, "::::::::::::::*:"),
	(0,     0,     0,     ':',     5,     0, ":::B::::::::::*:"),
	(0,     0,     1,     'B',     7,     0, ":::B::::::::::*:"),
	(0,     0,     1,     'W',     7,     0, ":::B:::B::::::*:"),
	(0,     0,     1,     '*',     7,     0, ":::B:::W::::::*:"),
	(0,     0,     0,     '*',     12,     0, ":::B:::B::::::*:"),
	(0,     1,     0,     '*',     1,     0, ":::B:::B::::::*:"),
	(0,     0,     0,     'B',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     3,     0, "::::W:::::::::::"),
	(0,     0,     1,     'W',     4,     0, ":::BW:::::::::::"),
	(0,     0,     0,     ':',     0,     0, ":::BW:::::::::::"),
	(0,     0,     0,     'W',     2,     0, ":::BW:::::::::::"),
	(0,     0,     1,     'W',     12,     0, ":::BW:::::::::::"),
	(0,     0,     0,     ':',     6,     0, ":::BW:::::::W:::"),
	(0,     0,     1,     '*',     13,     0, ":::BW:::::::W:::"),
	(0,     1,     1,     'W',     10,     0, ":::BW:::::::W*::"),
	(0,     0,     0,     '*',     10,     0, "::::::::::W:::::"),
	(0,     0,     0,     ':',     14,     0, "::::::::::W:::::"),
	(0,     0,     0,     'B',     10,     0, "::::::::::W:::::"),
	(0,     0,     1,     '*',     1,     0, "::::::::::W:::::"),
	(0,     0,     1,     'W',     10,     0, ":*::::::::W:::::"),
	(0,     0,     0,     '*',     2,     0, ":*::::::::W:::::"),
	(0,     0,     1,     'B',     2,     0, ":*::::::::W:::::"),
	(0,     0,     1,     ':',     11,     0, ":*B:::::::W:::::"),
	(0,     0,     0,     'W',     10,     0, ":*B:::::::W:::::"),
	(0,     0,     1,     ':',     3,     0, ":*B:::::::W:::::"),
	(0,     0,     1,     ':',     9,     0, ":*B:::::::W:::::"),
	(0,     0,     0,     'W',     7,     0, ":*B:::::::W:::::"),
	(0,     0,     1,     '*',     11,     0, ":*B:::::::W:::::"),
	(0,     0,     1,     'W',     5,     0, ":*B:::::::W*::::"),
	(0,     1,     1,     'B',     10,     0, ":*B::W::::W*::::"),
	(0,     0,     0,     'W',     8,     0, "::::::::::B:::::"),
	(0,     0,     0,     ':',     3,     0, "::::::::::B:::::"),
	(0,     0,     0,     '*',     1,     0, "::::::::::B:::::"),
	(0,     0,     1,     '*',     1,     0, "::::::::::B:::::"),
	(0,     0,     1,     ':',     1,     0, ":*::::::::B:::::"),
	(0,     0,     0,     'B',     3,     0, ":*::::::::B:::::"),
	(0,     0,     1,     'W',     13,     0, ":*::::::::B:::::"),
	(0,     0,     0,     'W',     0,     0, ":*::::::::B::W::"),
	(0,     1,     0,     'W',     13,     0, ":*::::::::B::W::"),
	(0,     0,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     2,     0, "B:::::::::::::::"),
	(0,     0,     0,     'W',     15,     0, "B:::::::::::::::"),
	(0,     1,     0,     ':',     12,     0, "B:::::::::::::::"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     0,     0, ":::::W::::::::::"),
	(0,     0,     1,     'B',     0,     0, "*::::W::::::::::"),
	(0,     0,     0,     ':',     5,     0, "B::::W::::::::::"),
	(0,     0,     0,     'B',     5,     0, "B::::W::::::::::"),
	(0,     0,     1,     'W',     13,     0, "B::::W::::::::::"),
	(0,     0,     1,     '*',     5,     0, "B::::W:::::::W::"),
	(0,     0,     1,     ':',     1,     0, "B::::B:::::::W::"),
	(0,     0,     0,     '*',     8,     0, "B::::B:::::::W::"),
	(0,     0,     1,     'W',     9,     0, "B::::B:::::::W::"),
	(0,     0,     1,     ':',     8,     0, "B::::B:::W:::W::"),
	(0,     0,     1,     'W',     5,     0, "B::::B:::W:::W::"),
	(1,     0,     1,     'B',     14,     0, "B::::W:::W:::W::"),
	(0,     0,     0,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     6,     0, ":::::::::::::W::"),
	(0,     0,     0,     '*',     13,     0, ":::::::::::::W::"),
	(0,     0,     0,     'W',     1,     0, ":::::::::::::W::"),
	(0,     1,     0,     'B',     0,     0, ":::::::::::::W::"),
	(0,     0,     0,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     11,     0, ":::::::::::B::::"),
	(0,     0,     1,     'B',     1,     0, ":::::::::::B::::"),
	(0,     0,     1,     'W',     14,     0, ":B:::::::::B::::"),
	(0,     0,     0,     ':',     12,     0, ":B:::::::::B::W:"),
	(0,     0,     0,     ':',     3,     0, ":B:::::::::B::W:"),
	(0,     0,     0,     'W',     0,     0, ":B:::::::::B::W:"),
	(0,     0,     0,     ':',     1,     0, ":B:::::::::B::W:"),
	(0,     0,     1,     'W',     13,     0, ":B:::::::::B::W:"),
	(0,     0,     1,     '*',     12,     0, ":B:::::::::B:WW:"),
	(0,     0,     0,     'W',     15,     0, ":B:::::::::B*WW:"),
	(0,     0,     0,     ':',     2,     0, ":B:::::::::B*WW:"),
	(0,     0,     0,     'W',     11,     0, ":B:::::::::B*WW:"),
	(0,     1,     0,     'W',     3,     0, ":B:::::::::B*WW:"),
	(0,     0,     1,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     13,     0, ":::::::::*::::::"),
	(0,     0,     1,     'W',     3,     0, ":::::::::*:::*::"),
	(0,     0,     1,     'W',     14,     0, ":::W:::::*:::*::"),
	(0,     0,     1,     ':',     4,     0, ":::W:::::*:::*W:"),
	(0,     0,     1,     ':',     6,     0, ":::W:::::*:::*W:"),
	(0,     0,     0,     '*',     12,     0, ":::W:::::*:::*W:"),
	(0,     0,     0,     '*',     12,     0, ":::W:::::*:::*W:"),
	(0,     0,     1,     'W',     13,     0, ":::W:::::*:::*W:"),
	(0,     0,     1,     ':',     6,     0, ":::W:::::*:::WW:"),
	(0,     0,     1,     'W',     12,     0, ":::W:::::*:::WW:"),
	(0,     0,     0,     'B',     1,     0, ":::W:::::*::WWW:"),
	(0,     0,     0,     'B',     0,     0, ":::W:::::*::WWW:"),
	(0,     0,     1,     'W',     7,     0, ":::W:::::*::WWW:"),
	(0,     0,     1,     ':',     5,     0, ":::W:::W:*::WWW:"),
	(0,     0,     0,     ':',     14,     0, ":::W:::W:*::WWW:"),
	(0,     0,     1,     'B',     7,     0, ":::W:::W:*::WWW:"),
	(0,     0,     0,     'B',     11,     0, ":::W:::B:*::WWW:"),
	(0,     0,     0,     'W',     8,     0, ":::W:::B:*::WWW:"),
	(0,     0,     1,     '*',     4,     0, ":::W:::B:*::WWW:"),
	(0,     0,     0,     '*',     3,     0, ":::W*::B:*::WWW:"),
	(0,     0,     0,     '*',     0,     0, ":::W*::B:*::WWW:"),
	(0,     0,     1,     'B',     2,     0, ":::W*::B:*::WWW:"),
	(0,     1,     1,     '*',     1,     0, "::BW*::B:*::WWW:"),
	(0,     0,     0,     '*',     15,     0, ":*::::::::::::::"),
	(0,     0,     0,     'B',     14,     0, ":*::::::::::::::"),
	(0,     0,     0,     'B',     5,     0, ":*::::::::::::::"),
	(0,     0,     0,     '*',     6,     0, ":*::::::::::::::"),
	(0,     1,     1,     'B',     12,     0, ":*::::::::::::::"),
	(0,     0,     0,     'B',     15,     0, "::::::::::::B:::"),
	(0,     0,     0,     'W',     12,     0, "::::::::::::B:::"),
	(0,     0,     1,     'B',     0,     0, "::::::::::::B:::"),
	(0,     0,     0,     'B',     2,     0, "B:::::::::::B:::"),
	(0,     0,     0,     '*',     10,     0, "B:::::::::::B:::"),
	(0,     0,     0,     'W',     14,     0, "B:::::::::::B:::"),
	(0,     0,     1,     '*',     13,     0, "B:::::::::::B:::"),
	(0,     1,     0,     ':',     13,     0, "B:::::::::::B*::"),
	(0,     0,     1,     'B',     15,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     7,     0, ":::::::::::::::B"),
	(0,     0,     0,     ':',     14,     0, ":::::::*:::::::B"),
	(0,     0,     1,     'B',     14,     0, ":::::::*:::::::B"),
	(0,     0,     1,     'W',     10,     0, ":::::::*::::::BB"),
	(0,     0,     0,     ':',     9,     0, ":::::::*::W:::BB"),
	(0,     0,     1,     'B',     14,     0, ":::::::*::W:::BB"),
	(0,     0,     1,     ':',     2,     0, ":::::::*::W:::BB"),
	(0,     0,     0,     '*',     2,     0, ":::::::*::W:::BB"),
	(0,     0,     1,     ':',     6,     0, ":::::::*::W:::BB"),
	(0,     0,     1,     'W',     2,     0, ":::::::*::W:::BB"),
	(0,     0,     1,     '*',     2,     0, "::W::::*::W:::BB"),
	(0,     0,     1,     ':',     11,     0, "::B::::*::W:::BB"),
	(0,     0,     0,     'B',     0,     0, "::B::::*::W:::BB"),
	(0,     0,     0,     '*',     10,     0, "::B::::*::W:::BB"),
	(0,     0,     0,     ':',     5,     0, "::B::::*::W:::BB"),
	(0,     0,     0,     'W',     11,     0, "::B::::*::W:::BB"),
	(0,     0,     0,     'W',     11,     0, "::B::::*::W:::BB"),
	(0,     0,     0,     'B',     2,     0, "::B::::*::W:::BB"),
	(0,     1,     1,     '*',     13,     0, "::B::::*::W:::BB"),
	(0,     0,     0,     'W',     2,     0, ":::::::::::::*::"),
	(0,     0,     0,     'W',     5,     0, ":::::::::::::*::"),
	(0,     0,     1,     '*',     6,     0, ":::::::::::::*::"),
	(0,     0,     1,     'W',     1,     0, "::::::*::::::*::"),
	(0,     0,     1,     'W',     9,     0, ":W::::*::::::*::"),
	(0,     0,     1,     ':',     5,     0, ":W::::*::W:::*::"),
	(0,     1,     0,     'W',     7,     0, ":W::::*::W:::*::"),
	(0,     0,     1,     'B',     4,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     14,     0, "::::B:::::::::::"),
	(0,     0,     1,     'W',     6,     0, "::::::::::::::W:"),
	(0,     0,     0,     ':',     6,     0, "::::::W:::::::W:"),
	(0,     0,     0,     '*',     5,     0, "::::::W:::::::W:"),
	(0,     0,     1,     '*',     15,     0, "::::::W:::::::W:"),
	(0,     0,     1,     'B',     3,     0, "::::::W:::::::W*"),
	(0,     1,     0,     '*',     11,     0, ":::B::W:::::::W*"),
	(0,     0,     0,     '*',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     13,     0, "::::::::::*:::::"),
	(0,     0,     1,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     0,     0, "W:::::::::::::::"),
	(0,     0,     0,     'B',     5,     0, "W:::::::::::::::"),
	(0,     1,     0,     '*',     15,     0, "W:::::::::::::::"),
	(0,     0,     1,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     4,     0, ":::::::::*::::::"),
	(0,     0,     0,     '*',     5,     0, ":::::::::*::::::"),
	(0,     0,     1,     ':',     6,     0, ":::::::::*::::::"),
	(0,     0,     0,     'W',     3,     0, ":::::::::*::::::"),
	(0,     0,     0,     'W',     12,     0, ":::::::::*::::::"),
	(0,     1,     1,     '*',     5,     0, ":::::::::*::::::"),
	(0,     1,     1,     ':',     10,     0, ":::::*::::::::::"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     11,     0, ":::::::::*::::::"),
	(0,     0,     1,     '*',     8,     0, ":::::::::*::::::"),
	(0,     0,     1,     '*',     9,     0, "::::::::**::::::"),
	(0,     0,     0,     ':',     3,     0, "::::::::*:::::::"),
	(0,     0,     0,     ':',     12,     0, "::::::::*:::::::"),
	(0,     0,     1,     'W',     15,     0, "::::::::*:::::::"),
	(0,     0,     0,     ':',     4,     0, "::::::::*::::::W"),
	(0,     0,     1,     '*',     14,     0, "::::::::*::::::W"),
	(0,     0,     1,     ':',     5,     0, "::::::::*:::::*W"),
	(0,     0,     0,     'W',     5,     0, "::::::::*:::::*W"),
	(0,     0,     0,     '*',     6,     0, "::::::::*:::::*W"),
	(0,     0,     1,     ':',     1,     0, "::::::::*:::::*W"),
	(0,     1,     1,     'W',     12,     0, "::::::::*:::::*W"),
	(0,     0,     0,     '*',     11,     0, "::::::::::::W:::"),
	(0,     0,     1,     'W',     13,     0, "::::::::::::W:::"),
	(0,     0,     0,     ':',     15,     0, "::::::::::::WW::"),
	(0,     0,     0,     'B',     12,     0, "::::::::::::WW::"),
	(0,     0,     1,     'B',     13,     0, "::::::::::::WW::"),
	(0,     0,     1,     'B',     13,     0, "::::::::::::WB::"),
	(0,     0,     0,     '*',     2,     0, "::::::::::::WB::"),
	(0,     0,     0,     '*',     8,     0, "::::::::::::WB::"),
	(0,     0,     0,     ':',     2,     0, "::::::::::::WB::"),
	(0,     0,     0,     'B',     14,     0, "::::::::::::WB::"),
	(0,     0,     0,     '*',     7,     0, "::::::::::::WB::"),
	(0,     1,     0,     'W',     8,     0, "::::::::::::WB::"),
	(0,     0,     0,     'B',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     1,     1, "::::::::::::::::"),
	(0,     1,     0,     'W',     1,     0, ":B::::::::::::::"),
	(0,     0,     1,     '*',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     14,     0, ":::::::::::*::::"),
	(0,     0,     0,     'W',     12,     0, ":::::::::::*::::"),
	(0,     0,     0,     ':',     15,     0, ":::::::::::*::::"),
	(0,     0,     0,     'W',     7,     0, ":::::::::::*::::"),
	(0,     0,     0,     '*',     13,     0, ":::::::::::*::::"),
	(0,     0,     0,     'W',     8,     0, ":::::::::::*::::"),
	(0,     0,     1,     'B',     11,     0, ":::::::::::*::::"),
	(0,     0,     1,     'W',     13,     0, ":::::::::::B::::"),
	(0,     0,     1,     'W',     0,     0, ":::::::::::B:W::"),
	(0,     1,     1,     'B',     10,     0, "W::::::::::B:W::"),
	(0,     0,     0,     'B',     1,     0, "::::::::::B:::::"),
	(0,     1,     1,     'B',     6,     0, "::::::::::B:::::"),
	(0,     0,     1,     'B',     0,     0, "::::::B:::::::::"),
	(0,     0,     1,     'W',     14,     0, "B:::::B:::::::::"),
	(0,     0,     0,     'B',     2,     0, "B:::::B:::::::W:"),
	(0,     0,     0,     'W',     4,     0, "B:::::B:::::::W:"),
	(0,     0,     1,     'B',     15,     0, "B:::::B:::::::W:"),
	(0,     0,     0,     'W',     15,     0, "B:::::B:::::::WB"),
	(0,     1,     0,     'W',     10,     0, "B:::::B:::::::WB"),
	(0,     0,     0,     'B',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     12,     0, "B:::::::::::::::"),
	(0,     0,     1,     'B',     8,     0, "B:::::::::::*:::"),
	(0,     0,     1,     'W',     9,     0, "B:::::::B:::*:::"),
	(0,     0,     1,     ':',     3,     0, "B:::::::BW::*:::"),
	(0,     0,     1,     'B',     0,     0, "B:::::::BW::*:::"),
	(0,     1,     1,     ':',     10,     0, "B:::::::BW::*:::"),
	(0,     0,     0,     '*',     6,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     15,     0, "::::::::::*:::::"),
	(0,     0,     1,     '*',     6,     0, "::::::::::*:::::"),
	(0,     0,     1,     '*',     4,     0, "::::::*:::*:::::"),
	(0,     0,     1,     '*',     12,     0, "::::*:*:::*:::::"),
	(0,     0,     1,     'B',     2,     0, "::::*:*:::*:*:::"),
	(0,     1,     0,     '*',     3,     0, "::B:*:*:::*:*:::"),
	(0,     0,     1,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     12,     0, ":::::::::::::::W"),
	(0,     0,     0,     'B',     3,     0, ":::::::::::::::W"),
	(0,     0,     1,     'W',     12,     0, ":::::::::::::::W"),
	(0,     0,     0,     'B',     14,     0, "::::::::::::W::W"),
	(0,     0,     0,     'B',     10,     0, "::::::::::::W::W"),
	(0,     0,     0,     'B',     4,     0, "::::::::::::W::W"),
	(0,     0,     1,     '*',     6,     0, "::::::::::::W::W"),
	(0,     1,     1,     'W',     4,     0, "::::::*:::::W::W"),
	(0,     0,     1,     '*',     9,     0, "::::W:::::::::::"),
	(0,     0,     1,     'B',     6,     0, "::::W::::*::::::"),
	(0,     0,     1,     ':',     5,     0, "::::W:B::*::::::"),
	(0,     0,     1,     'B',     5,     0, "::::W:B::*::::::"),
	(0,     0,     1,     'B',     11,     0, "::::WBB::*::::::"),
	(0,     0,     1,     '*',     5,     0, "::::WBB::*:B::::"),
	(0,     0,     1,     ':',     7,     0, "::::WWB::*:B::::"),
	(0,     0,     1,     'B',     14,     0, "::::WWB::*:B::::"),
	(0,     0,     0,     ':',     12,     0, "::::WWB::*:B::B:"),
	(0,     0,     0,     'B',     5,     0, "::::WWB::*:B::B:"),
	(0,     0,     0,     'W',     14,     0, "::::WWB::*:B::B:"),
	(0,     0,     0,     ':',     11,     0, "::::WWB::*:B::B:"),
	(0,     1,     1,     '*',     14,     0, "::::WWB::*:B::B:"),
	(0,     0,     0,     'B',     1,     0, "::::::::::::::*:"),
	(0,     0,     1,     'B',     6,     0, "::::::::::::::*:"),
	(0,     0,     1,     'B',     13,     0, "::::::B:::::::*:"),
	(0,     0,     0,     'W',     1,     0, "::::::B::::::B*:"),
	(0,     0,     0,     '*',     15,     0, "::::::B::::::B*:"),
	(0,     0,     1,     ':',     13,     0, "::::::B::::::B*:"),
	(0,     0,     1,     'W',     14,     0, "::::::B::::::B*:"),
	(0,     0,     1,     'B',     4,     0, "::::::B::::::BW:"),
	(0,     1,     0,     '*',     13,     0, "::::B:B::::::BW:"),
	(0,     0,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     15,     0, ":::::::::::*::::"),
	(0,     0,     1,     'B',     3,     0, ":::::::::::*:::W"),
	(0,     0,     0,     'W',     14,     0, ":::B:::::::*:::W"),
	(0,     1,     0,     ':',     0,     0, ":::B:::::::*:::W"),
	(0,     1,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     1,     0, "::::::W:::::::::"),
	(0,     0,     0,     ':',     14,     0, "::::::W:::::::::"),
	(0,     0,     0,     'B',     4,     0, "::::::W:::::::::"),
	(0,     0,     1,     'W',     0,     0, "::::::W:::::::::"),
	(0,     0,     1,     '*',     8,     0, "W:::::W:::::::::"),
	(0,     0,     1,     '*',     2,     0, "W:::::W:*:::::::"),
	(0,     0,     1,     'W',     7,     0, "W:*:::W:*:::::::"),
	(0,     0,     1,     '*',     3,     0, "W:*:::WW*:::::::"),
	(0,     0,     0,     '*',     4,     0, "W:**::WW*:::::::"),
	(0,     0,     0,     'W',     15,     0, "W:**::WW*:::::::"),
	(0,     0,     1,     'B',     8,     0, "W:**::WW*:::::::"),
	(0,     0,     1,     ':',     7,     0, "W:**::WWB:::::::"),
	(0,     0,     1,     'W',     15,     0, "W:**::WWB:::::::"),
	(0,     0,     1,     'B',     2,     0, "W:**::WWB::::::W"),
	(0,     0,     0,     'B',     4,     0, "W:B*::WWB::::::W"),
	(0,     0,     1,     'B',     0,     0, "W:B*::WWB::::::W"),
	(0,     0,     0,     'W',     2,     0, "B:B*::WWB::::::W"),
	(0,     0,     0,     ':',     1,     0, "B:B*::WWB::::::W"),
	(0,     0,     1,     '*',     2,     0, "B:B*::WWB::::::W"),
	(0,     0,     0,     '*',     7,     0, "B:W*::WWB::::::W"),
	(0,     0,     1,     'B',     13,     0, "B:W*::WWB::::::W"),
	(0,     0,     1,     'W',     3,     0, "B:W*::WWB::::B:W"),
	(0,     0,     0,     'W',     5,     0, "B:WW::WWB::::B:W"),
	(0,     0,     0,     'B',     15,     0, "B:WW::WWB::::B:W"),
	(0,     1,     1,     'W',     13,     0, "B:WW::WWB::::B:W"),
	(0,     0,     1,     '*',     10,     0, ":::::::::::::W::"),
	(0,     0,     0,     ':',     2,     0, "::::::::::*::W::"),
	(0,     0,     1,     '*',     11,     0, "::::::::::*::W::"),
	(0,     0,     0,     ':',     8,     0, "::::::::::**:W::"),
	(0,     0,     1,     'B',     13,     0, "::::::::::**:W::"),
	(0,     0,     0,     'B',     9,     0, "::::::::::**:B::"),
	(0,     0,     0,     'B',     11,     0, "::::::::::**:B::"),
	(0,     1,     1,     'B',     14,     0, "::::::::::**:B::"),
	(0,     0,     0,     '*',     13,     0, "::::::::::::::B:"),
	(0,     1,     0,     ':',     12,     0, "::::::::::::::B:"),
	(0,     0,     1,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     12,     0, "::::::::::::::W:"),
	(0,     0,     0,     '*',     14,     0, "::::::::::::*:W:"),
	(0,     0,     1,     '*',     0,     0, "::::::::::::*:W:"),
	(0,     1,     1,     'B',     8,     0, "*:::::::::::*:W:"),
	(0,     0,     1,     'B',     15,     0, "::::::::B:::::::"),
	(0,     0,     1,     ':',     7,     0, "::::::::B::::::B"),
	(0,     1,     0,     ':',     6,     0, "::::::::B::::::B"),
	(0,     0,     1,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     15,     0, "W:::::::::::::::"),
	(0,     0,     1,     '*',     6,     0, "W:::::::::::::::"),
	(0,     0,     0,     '*',     9,     0, "W:::::*:::::::::"),
	(0,     1,     1,     'W',     13,     0, "W:::::*:::::::::"),
	(0,     1,     1,     '*',     14,     0, ":::::::::::::W::"),
	(0,     1,     1,     '*',     15,     0, "::::::::::::::*:"),
	(0,     0,     1,     'W',     14,     0, ":::::::::::::::*"),
	(0,     0,     1,     'B',     10,     0, "::::::::::::::W*"),
	(0,     1,     1,     'B',     7,     0, "::::::::::B:::W*"),
	(0,     0,     0,     ':',     9,     0, ":::::::B::::::::"),
	(0,     0,     1,     'W',     1,     0, ":::::::B::::::::"),
	(0,     0,     1,     ':',     10,     0, ":W:::::B::::::::"),
	(0,     0,     0,     'B',     9,     0, ":W:::::B::::::::"),
	(0,     0,     0,     'B',     12,     0, ":W:::::B::::::::"),
	(0,     0,     0,     '*',     1,     0, ":W:::::B::::::::"),
	(0,     0,     1,     ':',     13,     0, ":W:::::B::::::::"),
	(0,     0,     1,     ':',     11,     0, ":W:::::B::::::::"),
	(0,     1,     1,     '*',     12,     0, ":W:::::B::::::::"),
	(0,     0,     1,     ':',     4,     0, "::::::::::::*:::"),
	(0,     0,     1,     ':',     9,     0, "::::::::::::*:::"),
	(0,     1,     0,     ':',     6,     0, "::::::::::::*:::"),
	(0,     0,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     10,     0, "::::::::::*:::::"),
	(0,     0,     1,     'B',     4,     0, "::::::::::*:::::"),
	(0,     1,     1,     'B',     3,     0, "::::B:::::*:::::"),
	(0,     0,     1,     '*',     4,     0, ":::B::::::::::::"),
	(0,     0,     0,     ':',     12,     0, ":::B*:::::::::::"),
	(0,     0,     1,     'B',     6,     0, ":::B*:::::::::::"),
	(0,     0,     1,     ':',     1,     0, ":::B*:B:::::::::"),
	(0,     0,     1,     'W',     3,     0, ":::B*:B:::::::::"),
	(0,     0,     0,     'B',     13,     0, ":::W*:B:::::::::"),
	(0,     0,     0,     ':',     7,     0, ":::W*:B:::::::::"),
	(0,     0,     1,     '*',     4,     0, ":::W*:B:::::::::"),
	(0,     0,     0,     '*',     13,     0, ":::W::B:::::::::"),
	(0,     0,     0,     'W',     10,     0, ":::W::B:::::::::"),
	(0,     0,     0,     'W',     15,     0, ":::W::B:::::::::"),
	(0,     0,     0,     '*',     9,     0, ":::W::B:::::::::"),
	(0,     0,     1,     'W',     12,     0, ":::W::B:::::::::"),
	(0,     0,     1,     'B',     1,     0, ":::W::B:::::W:::"),
	(0,     0,     0,     'W',     13,     0, ":B:W::B:::::W:::"),
	(0,     0,     0,     'W',     1,     0, ":B:W::B:::::W:::"),
	(0,     0,     0,     'W',     0,     0, ":B:W::B:::::W:::"),
	(0,     1,     1,     ':',     7,     0, ":B:W::B:::::W:::"),
	(0,     0,     1,     '*',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     8,     0, "::::::::::::*:::"),
	(0,     0,     1,     ':',     0,     0, "::::::::B:::*:::"),
	(0,     0,     0,     'B',     6,     0, "::::::::B:::*:::"),
	(0,     0,     1,     'W',     5,     0, "::::::::B:::*:::"),
	(0,     0,     0,     'W',     12,     0, ":::::W::B:::*:::"),
	(0,     0,     0,     'B',     5,     0, ":::::W::B:::*:::"),
	(0,     0,     0,     '*',     5,     0, ":::::W::B:::*:::"),
	(0,     1,     0,     '*',     15,     0, ":::::W::B:::*:::"),
	(0,     0,     0,     '*',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     5,     0, "::::::::::::W:::"),
	(0,     0,     1,     'B',     1,     0, "::::::::::::W:::"),
	(0,     0,     0,     ':',     11,     0, ":B::::::::::W:::"),
	(0,     0,     0,     '*',     5,     0, ":B::::::::::W:::"),
	(0,     0,     0,     ':',     7,     0, ":B::::::::::W:::"),
	(0,     0,     0,     'B',     4,     0, ":B::::::::::W:::"),
	(0,     0,     0,     'B',     2,     0, ":B::::::::::W:::"),
	(0,     0,     1,     'W',     10,     0, ":B::::::::::W:::"),
	(0,     1,     0,     ':',     8,     0, ":B::::::::W:W:::"),
	(0,     1,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     15,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     3,     0, "::::::W:::::::::"),
	(0,     0,     0,     'W',     10,     0, ":::B::W:::::::::"),
	(0,     0,     1,     '*',     14,     0, ":::B::W:::::::::"),
	(0,     0,     1,     '*',     14,     0, ":::B::W:::::::*:"),
	(0,     1,     1,     '*',     1,     0, ":::B::W:::::::::"),
	(0,     0,     0,     'W',     8,     0, ":*::::::::::::::"),
	(0,     0,     1,     'W',     11,     0, ":*::::::::::::::"),
	(0,     0,     0,     'B',     1,     0, ":*:::::::::W::::"),
	(0,     0,     0,     '*',     7,     0, ":*:::::::::W::::"),
	(0,     0,     1,     'B',     11,     0, ":*:::::::::W::::"),
	(0,     1,     1,     ':',     2,     0, ":*:::::::::B::::"),
	(0,     1,     1,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     6,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     1,     0, "::::::::::::::B:"),
	(0,     0,     0,     '*',     12,     0, "::::::::::::::B:"),
	(0,     0,     1,     '*',     10,     0, "::::::::::::::B:"),
	(0,     0,     1,     ':',     9,     0, "::::::::::*:::B:"),
	(0,     0,     0,     ':',     9,     0, "::::::::::*:::B:"),
	(0,     0,     0,     'B',     9,     0, "::::::::::*:::B:"),
	(0,     0,     0,     'B',     9,     0, "::::::::::*:::B:"),
	(0,     0,     1,     '*',     13,     0, "::::::::::*:::B:"),
	(0,     1,     1,     ':',     9,     0, "::::::::::*::*B:"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     14,     0, "*:::::::::::::::"),
	(0,     1,     0,     ':',     4,     0, "*:::::::::::::*:"),
	(0,     0,     0,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     6,     0, "::::::::B:::::::"),
	(0,     0,     1,     '*',     10,     0, "::::::::B:::::::"),
	(0,     0,     1,     ':',     5,     0, "::::::::B:*:::::"),
	(0,     0,     1,     ':',     12,     0, "::::::::B:*:::::"),
	(0,     0,     1,     '*',     13,     0, "::::::::B:*:::::"),
	(0,     0,     1,     ':',     12,     0, "::::::::B:*::*::"),
	(0,     0,     0,     '*',     0,     0, "::::::::B:*::*::"),
	(0,     0,     0,     'W',     14,     0, "::::::::B:*::*::"),
	(0,     0,     0,     '*',     0,     0, "::::::::B:*::*::"),
	(0,     1,     1,     '*',     3,     0, "::::::::B:*::*::"),
	(0,     1,     0,     'B',     14,     0, ":::*::::::::::::"),
	(0,     0,     0,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     4,     0, "*:::::::::::::::"),
	(0,     0,     0,     'W',     15,     0, "*:::::::::::::::"),
	(0,     0,     0,     'W',     1,     0, "*:::::::::::::::"),
	(0,     0,     1,     'B',     15,     0, "*:::::::::::::::"),
	(0,     1,     0,     'B',     12,     0, "*::::::::::::::B"),
	(0,     0,     1,     ':',     1,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     3,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     13,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     3,     0, ":::::*::::::::::"),
	(0,     0,     1,     'B',     1,     0, ":::::*::::::::::"),
	(0,     0,     1,     'W',     7,     0, ":B:::*::::::::::"),
	(0,     0,     0,     'B',     6,     0, ":B:::*:W::::::::"),
	(0,     0,     1,     ':',     12,     0, ":B:::*:W::::::::"),
	(0,     0,     1,     ':',     5,     0, ":B:::*:W::::::::"),
	(0,     1,     0,     ':',     11,     0, ":B:::*:W::::::::"),
	(0,     1,     0,     '*',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     5,     0, ":B::::::::::::::"),
	(0,     0,     0,     'W',     12,     0, ":B::::::::::::::"),
	(0,     1,     0,     '*',     2,     0, ":B::::::::::::::"),
	(0,     0,     1,     '*',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     4,     0, ":::::::::::*::::"),
	(0,     0,     1,     'W',     1,     0, ":::::::::::*::::"),
	(0,     0,     1,     ':',     8,     0, ":W:::::::::*::::"),
	(0,     0,     0,     'B',     7,     0, ":W:::::::::*::::"),
	(0,     0,     0,     'W',     3,     0, ":W:::::::::*::::"),
	(0,     0,     1,     'W',     15,     0, ":W:::::::::*::::"),
	(0,     0,     0,     'W',     3,     0, ":W:::::::::*:::W"),
	(0,     0,     1,     '*',     5,     0, ":W:::::::::*:::W"),
	(0,     0,     0,     'B',     12,     0, ":W:::*:::::*:::W"),
	(0,     1,     0,     'B',     3,     0, ":W:::*:::::*:::W"),
	(0,     0,     0,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     11,     0, ":::::::::::::B::"),
	(0,     0,     1,     '*',     15,     0, ":::::::::::::B::"),
	(0,     1,     0,     '*',     2,     0, ":::::::::::::B:*"),
	(0,     0,     1,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     5,     0, ":::::::::B::::::"),
	(0,     0,     0,     '*',     4,     0, ":::::::::B::::::"),
	(0,     0,     1,     ':',     12,     0, ":::::::::B::::::"),
	(0,     1,     0,     'B',     0,     0, ":::::::::B::::::"),
	(0,     0,     0,     ':',     6,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     7,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     9,     0, "::::::::::::::B:"),
	(0,     0,     0,     '*',     10,     0, ":::::::::B::::B:"),
	(0,     0,     0,     'W',     5,     0, ":::::::::B::::B:"),
	(0,     0,     0,     'B',     15,     0, ":::::::::B::::B:"),
	(0,     0,     1,     '*',     15,     0, ":::::::::B::::B:"),
	(0,     0,     0,     'W',     1,     0, ":::::::::B::::B*"),
	(0,     0,     0,     ':',     9,     0, ":::::::::B::::B*"),
	(0,     0,     1,     'B',     10,     0, ":::::::::B::::B*"),
	(0,     0,     0,     '*',     13,     0, ":::::::::BB:::B*"),
	(0,     0,     0,     'B',     14,     0, ":::::::::BB:::B*"),
	(0,     0,     0,     ':',     4,     0, ":::::::::BB:::B*"),
	(0,     0,     0,     'W',     10,     0, ":::::::::BB:::B*"),
	(0,     0,     1,     ':',     3,     0, ":::::::::BB:::B*"),
	(0,     0,     0,     ':',     12,     0, ":::::::::BB:::B*"),
	(0,     0,     1,     '*',     3,     0, ":::::::::BB:::B*"),
	(0,     0,     0,     'W',     13,     0, ":::*:::::BB:::B*"),
	(0,     0,     0,     ':',     8,     0, ":::*:::::BB:::B*"),
	(0,     0,     1,     ':',     5,     0, ":::*:::::BB:::B*"),
	(0,     0,     0,     '*',     15,     0, ":::*:::::BB:::B*"),
	(0,     0,     1,     ':',     3,     0, ":::*:::::BB:::B*"),
	(0,     0,     0,     'B',     15,     0, ":::*:::::BB:::B*"),
	(0,     0,     1,     ':',     2,     0, ":::*:::::BB:::B*"),
	(0,     0,     0,     'B',     2,     0, ":::*:::::BB:::B*"),
	(0,     1,     0,     'B',     0,     0, ":::*:::::BB:::B*"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     14,     0, "::::::*:::::::::"),
	(0,     0,     1,     'B',     10,     0, "::::::*:::::::::"),
	(0,     0,     0,     'B',     11,     0, "::::::*:::B:::::"),
	(0,     0,     0,     ':',     15,     0, "::::::*:::B:::::"),
	(0,     0,     0,     'W',     2,     0, "::::::*:::B:::::"),
	(0,     0,     0,     'W',     8,     0, "::::::*:::B:::::"),
	(0,     0,     0,     '*',     12,     0, "::::::*:::B:::::"),
	(0,     0,     1,     'B',     5,     0, "::::::*:::B:::::"),
	(0,     0,     1,     'W',     15,     0, ":::::B*:::B:::::"),
	(0,     0,     0,     '*',     4,     0, ":::::B*:::B::::W"),
	(0,     0,     0,     ':',     6,     0, ":::::B*:::B::::W"),
	(0,     0,     0,     '*',     0,     0, ":::::B*:::B::::W"),
	(0,     0,     0,     ':',     10,     0, ":::::B*:::B::::W"),
	(0,     0,     1,     'W',     7,     0, ":::::B*:::B::::W"),
	(0,     0,     1,     'W',     5,     0, ":::::B*W::B::::W"),
	(0,     0,     0,     '*',     5,     0, ":::::W*W::B::::W"),
	(0,     1,     1,     'W',     15,     0, ":::::W*W::B::::W"),
	(0,     0,     1,     'B',     9,     0, ":::::::::::::::W"),
	(0,     0,     1,     '*',     9,     0, ":::::::::B:::::W"),
	(0,     0,     1,     'B',     2,     0, ":::::::::W:::::W"),
	(0,     0,     0,     'W',     11,     0, "::B::::::W:::::W"),
	(0,     1,     1,     '*',     0,     0, "::B::::::W:::::W"),
	(0,     0,     0,     '*',     14,     0, "*:::::::::::::::"),
	(0,     1,     0,     '*',     11,     0, "*:::::::::::::::"),
	(0,     0,     1,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     6,     0, "::::::::::W:::::"),
	(0,     0,     0,     'W',     5,     0, "::::::B:::W:::::"),
	(0,     0,     1,     'B',     1,     0, "::::::B:::W:::::"),
	(0,     0,     0,     'B',     13,     0, ":B::::B:::W:::::"),
	(0,     0,     0,     'B',     9,     0, ":B::::B:::W:::::"),
	(0,     0,     1,     'W',     10,     0, ":B::::B:::W:::::"),
	(0,     0,     1,     'W',     13,     0, ":B::::B:::W:::::"),
	(0,     1,     1,     'B',     9,     0, ":B::::B:::W::W::"),
	(0,     0,     1,     'W',     14,     0, ":::::::::B::::::"),
	(0,     0,     0,     ':',     11,     0, ":::::::::B::::W:"),
	(0,     0,     0,     'W',     12,     0, ":::::::::B::::W:"),
	(0,     0,     1,     'W',     7,     0, ":::::::::B::::W:"),
	(0,     0,     0,     'W',     2,     0, ":::::::W:B::::W:"),
	(0,     0,     0,     'B',     0,     0, ":::::::W:B::::W:"),
	(0,     1,     0,     ':',     14,     0, ":::::::W:B::::W:"),
	(0,     0,     1,     'W',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     10,     0, ":::::::::::W::::"),
	(0,     0,     0,     '*',     3,     0, ":::::::::::W::::"),
	(0,     0,     0,     'B',     2,     0, ":::::::::::W::::"),
	(0,     0,     1,     '*',     11,     0, ":::::::::::W::::"),
	(0,     0,     0,     ':',     4,     0, ":::::::::::B::::"),
	(0,     0,     0,     '*',     12,     0, ":::::::::::B::::"),
	(0,     0,     0,     ':',     7,     0, ":::::::::::B::::"),
	(0,     0,     0,     'W',     13,     0, ":::::::::::B::::"),
	(0,     0,     0,     'B',     5,     0, ":::::::::::B::::"),
	(0,     0,     0,     'B',     6,     0, ":::::::::::B::::"),
	(0,     1,     1,     'W',     15,     0, ":::::::::::B::::"),
	(0,     0,     0,     'W',     9,     0, ":::::::::::::::W"),
	(0,     0,     0,     '*',     15,     0, ":::::::::::::::W"),
	(0,     0,     1,     'W',     15,     0, ":::::::::::::::W"),
	(0,     0,     0,     'W',     6,     0, ":::::::::::::::W"),
	(0,     0,     1,     '*',     2,     0, ":::::::::::::::W"),
	(0,     0,     0,     '*',     14,     0, "::*::::::::::::W"),
	(0,     0,     0,     'W',     13,     0, "::*::::::::::::W"),
	(0,     0,     0,     'B',     12,     0, "::*::::::::::::W"),
	(0,     0,     1,     '*',     7,     0, "::*::::::::::::W"),
	(0,     1,     0,     ':',     8,     0, "::*::::*:::::::W"),
	(0,     1,     0,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     2,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     11,     0, "::B:::::::::::::"),
	(0,     0,     1,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     7,     0, ":::::::W::::::::"),
	(0,     0,     1,     ':',     14,     0, ":::::::W::::::::"),
	(0,     1,     0,     '*',     12,     0, ":::::::W::::::::"),
	(0,     0,     1,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     15,     0, "::::W:::::::::::"),
	(0,     0,     1,     'W',     9,     0, "::::W::::::::::*"),
	(1,     1,     1,     ':',     2,     0, "::::W::::W:::::*"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     4,     0, ":::::::::B::::::"),
	(0,     0,     1,     'W',     10,     0, ":::::::::B::::::"),
	(0,     0,     1,     ':',     13,     0, ":::::::::BW:::::"),
	(0,     0,     0,     '*',     10,     0, ":::::::::BW:::::"),
	(0,     1,     1,     '*',     9,     0, ":::::::::BW:::::"),
	(0,     0,     1,     '*',     12,     0, ":::::::::*::::::"),
	(0,     0,     0,     'W',     12,     0, ":::::::::*::*:::"),
	(0,     0,     0,     ':',     11,     0, ":::::::::*::*:::"),
	(0,     0,     1,     ':',     7,     0, ":::::::::*::*:::"),
	(0,     0,     1,     'B',     12,     0, ":::::::::*::*:::"),
	(0,     0,     1,     'B',     0,     0, ":::::::::*::B:::"),
	(0,     0,     0,     'W',     10,     0, "B::::::::*::B:::"),
	(0,     0,     1,     '*',     7,     0, "B::::::::*::B:::"),
	(0,     0,     0,     ':',     1,     0, "B::::::*:*::B:::"),
	(0,     0,     1,     ':',     5,     0, "B::::::*:*::B:::"),
	(0,     0,     0,     ':',     5,     0, "B::::::*:*::B:::"),
	(0,     0,     0,     'B',     9,     0, "B::::::*:*::B:::"),
	(0,     0,     1,     '*',     13,     0, "B::::::*:*::B:::"),
	(0,     0,     1,     '*',     2,     0, "B::::::*:*::B*::"),
	(0,     0,     1,     'B',     0,     0, "B:*::::*:*::B*::"),
	(0,     1,     1,     '*',     6,     0, "B:*::::*:*::B*::"),
	(0,     0,     0,     '*',     0,     0, "::::::*:::::::::"),
	(0,     0,     0,     'B',     0,     0, "::::::*:::::::::"),
	(0,     0,     0,     'W',     12,     0, "::::::*:::::::::"),
	(0,     0,     0,     'W',     5,     0, "::::::*:::::::::"),
	(0,     0,     1,     'B',     10,     0, "::::::*:::::::::"),
	(0,     0,     1,     ':',     1,     0, "::::::*:::B:::::"),
	(0,     0,     1,     'B',     7,     0, "::::::*:::B:::::"),
	(0,     0,     0,     ':',     15,     0, "::::::*B::B:::::"),
	(0,     0,     0,     ':',     3,     0, "::::::*B::B:::::"),
	(0,     0,     0,     'W',     6,     0, "::::::*B::B:::::"),
	(0,     0,     1,     '*',     9,     0, "::::::*B::B:::::"),
	(0,     1,     1,     '*',     13,     0, "::::::*B:*B:::::"),
	(0,     0,     0,     'W',     1,     0, ":::::::::::::*::"),
	(0,     0,     0,     'B',     6,     0, ":::::::::::::*::"),
	(0,     0,     0,     '*',     4,     0, ":::::::::::::*::"),
	(0,     1,     1,     ':',     15,     0, ":::::::::::::*::"),
	(0,     0,     1,     ':',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     14,     0, "::*:::::::::::::"),
	(0,     0,     0,     ':',     11,     0, "::*:::::::::::::"),
	(0,     0,     0,     '*',     6,     0, "::*:::::::::::::"),
	(0,     0,     0,     ':',     10,     0, "::*:::::::::::::"),
	(0,     0,     0,     'W',     14,     0, "::*:::::::::::::"),
	(0,     0,     0,     'W',     9,     0, "::*:::::::::::::"),
	(0,     0,     0,     'B',     12,     0, "::*:::::::::::::"),
	(0,     0,     1,     'B',     15,     0, "::*:::::::::::::"),
	(0,     0,     1,     'B',     1,     0, "::*::::::::::::B"),
	(0,     0,     1,     'B',     10,     0, ":B*::::::::::::B"),
	(0,     0,     1,     'W',     15,     0, ":B*:::::::B::::B"),
	(0,     0,     1,     ':',     1,     0, ":B*:::::::B::::W"),
	(0,     0,     1,     'W',     9,     0, ":B*:::::::B::::W"),
	(0,     0,     1,     'B',     14,     0, ":B*::::::WB::::W"),
	(0,     1,     1,     ':',     4,     0, ":B*::::::WB:::BW"),
	(0,     1,     1,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     7,     0, ":::B::::::::::::"),
	(0,     0,     0,     'W',     6,     0, ":::B:::W::::::::"),
	(0,     0,     1,     'B',     6,     0, ":::B:::W::::::::"),
	(0,     0,     1,     ':',     2,     0, ":::B::BW::::::::"),
	(0,     0,     1,     '*',     8,     0, ":::B::BW::::::::"),
	(0,     0,     0,     ':',     5,     0, ":::B::BW*:::::::"),
	(0,     0,     0,     ':',     12,     0, ":::B::BW*:::::::"),
	(0,     0,     0,     '*',     12,     0, ":::B::BW*:::::::"),
	(0,     0,     0,     'B',     2,     0, ":::B::BW*:::::::"),
	(0,     0,     1,     ':',     8,     0, ":::B::BW*:::::::"),
	(0,     0,     0,     ':',     3,     0, ":::B::BW*:::::::"),
	(0,     0,     0,     'W',     9,     0, ":::B::BW*:::::::"),
	(0,     0,     0,     'W',     6,     0, ":::B::BW*:::::::"),
	(0,     0,     0,     'W',     2,     0, ":::B::BW*:::::::"),
	(0,     1,     0,     'W',     1,     0, ":::B::BW*:::::::"),
	(0,     0,     0,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     10,     0, ":B::::::::::::::"),
	(0,     0,     1,     ':',     5,     0, ":B::::::::::::::"),
	(0,     0,     0,     'W',     11,     0, ":B::::::::::::::"),
	(0,     0,     1,     'W',     9,     0, ":B::::::::::::::"),
	(0,     0,     0,     ':',     0,     0, ":B:::::::W::::::"),
	(0,     0,     1,     ':',     3,     0, ":B:::::::W::::::"),
	(0,     0,     1,     '*',     10,     0, ":B:::::::W::::::"),
	(0,     0,     0,     'B',     7,     0, ":B:::::::W*:::::"),
	(0,     0,     1,     ':',     4,     0, ":B:::::::W*:::::"),
	(0,     0,     1,     'B',     14,     0, ":B:::::::W*:::::"),
	(0,     0,     1,     ':',     0,     0, ":B:::::::W*:::B:"),
	(0,     1,     1,     '*',     13,     0, ":B:::::::W*:::B:"),
	(0,     0,     1,     '*',     1,     0, ":::::::::::::*::"),
	(0,     0,     1,     'W',     12,     0, ":*:::::::::::*::"),
	(0,     0,     0,     'W',     9,     0, ":*::::::::::W*::"),
	(0,     0,     0,     '*',     4,     0, ":*::::::::::W*::"),
	(0,     0,     1,     'B',     6,     0, ":*::::::::::W*::"),
	(0,     0,     0,     'B',     3,     0, ":*::::B:::::W*::"),
	(0,     0,     0,     '*',     10,     0, ":*::::B:::::W*::"),
	(0,     1,     1,     'W',     10,     0, ":*::::B:::::W*::"),
	(0,     0,     0,     'B',     12,     0, "::::::::::W:::::"),
	(0,     0,     0,     '*',     12,     0, "::::::::::W:::::"),
	(0,     0,     1,     '*',     0,     0, "::::::::::W:::::"),
	(0,     0,     0,     'W',     2,     0, "*:::::::::W:::::"),
	(0,     0,     0,     '*',     5,     0, "*:::::::::W:::::"),
	(0,     0,     0,     ':',     12,     0, "*:::::::::W:::::"),
	(0,     0,     0,     ':',     9,     0, "*:::::::::W:::::"),
	(0,     1,     0,     ':',     8,     0, "*:::::::::W:::::"),
	(0,     0,     0,     '*',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     7,     0, "W:::::::::::::::"),
	(0,     0,     0,     '*',     0,     0, "W:::::::::::::::"),
	(0,     0,     0,     ':',     15,     0, "W:::::::::::::::"),
	(0,     0,     1,     '*',     6,     0, "W:::::::::::::::"),
	(0,     1,     0,     'B',     9,     0, "W:::::*:::::::::"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     7,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     11,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     14,     0, ":::::::::::::::B"),
	(0,     0,     0,     'W',     9,     0, ":::::::::::::::B"),
	(0,     0,     1,     ':',     8,     0, ":::::::::::::::B"),
	(0,     0,     1,     'W',     2,     0, ":::::::::::::::B"),
	(0,     0,     0,     'W',     12,     0, "::W::::::::::::B"),
	(0,     0,     0,     'B',     4,     0, "::W::::::::::::B"),
	(0,     0,     0,     ':',     5,     0, "::W::::::::::::B"),
	(0,     0,     0,     'W',     8,     0, "::W::::::::::::B"),
	(0,     0,     0,     'W',     3,     0, "::W::::::::::::B"),
	(0,     0,     1,     'B',     10,     0, "::W::::::::::::B"),
	(0,     0,     0,     '*',     11,     0, "::W:::::::B::::B"),
	(0,     0,     0,     ':',     4,     0, "::W:::::::B::::B"),
	(0,     0,     1,     ':',     13,     0, "::W:::::::B::::B"),
	(0,     0,     0,     '*',     4,     0, "::W:::::::B::::B"),
	(0,     0,     0,     'B',     0,     0, "::W:::::::B::::B"),
	(0,     0,     1,     'W',     15,     0, "::W:::::::B::::B"),
	(0,     0,     0,     ':',     13,     0, "::W:::::::B::::W"),
	(0,     0,     1,     '*',     8,     0, "::W:::::::B::::W"),
	(0,     0,     1,     ':',     5,     0, "::W:::::*:B::::W"),
	(0,     0,     0,     '*',     1,     0, "::W:::::*:B::::W"),
	(0,     0,     1,     ':',     9,     0, "::W:::::*:B::::W"),
	(0,     0,     0,     ':',     3,     0, "::W:::::*:B::::W"),
	(0,     0,     1,     'B',     12,     0, "::W:::::*:B::::W"),
	(0,     1,     0,     ':',     5,     0, "::W:::::*:B:B::W"),
	(0,     0,     0,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     0, ":::::::::B::::::"),
	(0,     0,     1,     ':',     4,     0, ":::::::::B::::::"),
	(0,     0,     0,     ':',     1,     0, ":::::::::B::::::"),
	(0,     0,     1,     'W',     1,     0, ":::::::::B::::::"),
	(0,     0,     1,     'B',     4,     0, ":W:::::::B::::::"),
	(0,     0,     0,     'W',     1,     0, ":W::B::::B::::::"),
	(0,     0,     0,     ':',     7,     0, ":W::B::::B::::::"),
	(0,     0,     1,     '*',     4,     0, ":W::B::::B::::::"),
	(0,     0,     0,     '*',     10,     0, ":W::W::::B::::::"),
	(0,     0,     0,     'W',     2,     0, ":W::W::::B::::::"),
	(0,     0,     0,     'B',     2,     0, ":W::W::::B::::::"),
	(0,     0,     1,     'W',     11,     0, ":W::W::::B::::::"),
	(0,     0,     0,     ':',     11,     0, ":W::W::::B:W::::"),
	(0,     1,     0,     'W',     8,     0, ":W::W::::B:W::::"),
	(0,     0,     1,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     1,     0, ":::::::::::::W::"),
	(0,     1,     1,     '*',     1,     0, ":::::::::::::W::"),
	(0,     1,     1,     'W',     15,     0, ":*::::::::::::::"),
	(0,     0,     1,     'W',     4,     0, ":::::::::::::::W"),
	(0,     0,     1,     ':',     5,     0, "::::W::::::::::W"),
	(0,     0,     0,     'W',     9,     0, "::::W::::::::::W"),
	(0,     0,     0,     'W',     11,     0, "::::W::::::::::W"),
	(0,     0,     1,     ':',     11,     0, "::::W::::::::::W"),
	(0,     1,     0,     ':',     4,     0, "::::W::::::::::W"),
	(0,     0,     1,     ':',     5,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     4,     0, "::::::B:::::::::"),
	(0,     1,     0,     'B',     0,     0, "::::::B:::::::::"),
	(0,     0,     0,     'B',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     2,     0, "::::::::::::W:::"),
	(0,     1,     1,     ':',     4,     0, "::::::::::::W:::"),
	(0,     0,     0,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     15,     0, "::::::::B:::::::"),
	(0,     0,     0,     '*',     14,     0, "::::::::B:::::::"),
	(0,     0,     0,     'B',     5,     0, "::::::::B:::::::"),
	(0,     0,     1,     'W',     13,     0, "::::::::B:::::::"),
	(0,     0,     0,     ':',     7,     0, "::::::::B::::W::"),
	(0,     0,     0,     '*',     0,     0, "::::::::B::::W::"),
	(0,     1,     1,     'W',     7,     0, "::::::::B::::W::"),
	(0,     1,     1,     ':',     5,     0, ":::::::W::::::::"),
	(0,     0,     0,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     13,     0, ":::::::::B::::::"),
	(0,     1,     0,     'B',     2,     0, ":::::::::B:::W::"),
	(0,     0,     0,     'B',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     6,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     7,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     4,     0, ":::::::*::::::::"),
	(0,     0,     1,     '*',     10,     0, "::::B::*::::::::"),
	(0,     0,     1,     'W',     6,     0, "::::B::*::*:::::"),
	(0,     0,     1,     '*',     9,     0, "::::B:W*::*:::::"),
	(0,     0,     1,     'W',     3,     0, "::::B:W*:**:::::"),
	(0,     0,     1,     '*',     8,     0, ":::WB:W*:**:::::"),
	(0,     0,     0,     '*',     1,     0, ":::WB:W****:::::"),
	(0,     0,     1,     'B',     6,     0, ":::WB:W****:::::"),
	(0,     0,     0,     'W',     5,     0, ":::WB:B****:::::"),
	(0,     0,     1,     '*',     4,     0, ":::WB:B****:::::"),
	(0,     0,     0,     ':',     9,     0, ":::WW:B****:::::"),
	(0,     0,     1,     ':',     10,     0, ":::WW:B****:::::"),
	(0,     0,     1,     '*',     3,     0, ":::WW:B****:::::"),
	(0,     0,     1,     ':',     3,     0, ":::BW:B****:::::"),
	(0,     0,     0,     'W',     10,     0, ":::BW:B****:::::"),
	(0,     0,     0,     'B',     12,     0, ":::BW:B****:::::"),
	(0,     0,     0,     'B',     1,     0, ":::BW:B****:::::"),
	(0,     0,     0,     '*',     9,     0, ":::BW:B****:::::"),
	(0,     0,     0,     '*',     14,     0, ":::BW:B****:::::"),
	(0,     0,     1,     'B',     3,     0, ":::BW:B****:::::"),
	(0,     0,     1,     ':',     14,     0, ":::BW:B****:::::"),
	(0,     0,     0,     '*',     15,     0, ":::BW:B****:::::"),
	(0,     0,     0,     '*',     3,     0, ":::BW:B****:::::"),
	(0,     0,     0,     'B',     6,     0, ":::BW:B****:::::"),
	(0,     0,     0,     'W',     14,     0, ":::BW:B****:::::"),
	(0,     0,     1,     '*',     8,     0, ":::BW:B****:::::"),
	(0,     0,     1,     'B',     6,     0, ":::BW:B*:**:::::"),
	(0,     0,     1,     'B',     0,     0, ":::BW:B*:**:::::"),
	(0,     0,     0,     ':',     7,     0, "B::BW:B*:**:::::"),
	(0,     0,     0,     'B',     14,     0, "B::BW:B*:**:::::"),
	(0,     0,     1,     'W',     14,     0, "B::BW:B*:**:::::"),
	(0,     0,     0,     ':',     10,     0, "B::BW:B*:**:::W:"),
	(0,     0,     1,     'W',     14,     0, "B::BW:B*:**:::W:"),
	(0,     0,     0,     'B',     6,     0, "B::BW:B*:**:::W:"),
	(0,     0,     1,     '*',     15,     0, "B::BW:B*:**:::W:"),
	(0,     1,     1,     '*',     7,     0, "B::BW:B*:**:::W*"),
	(0,     0,     0,     'B',     4,     0, ":::::::*::::::::"),
	(0,     0,     0,     '*',     5,     0, ":::::::*::::::::"),
	(0,     0,     1,     ':',     11,     0, ":::::::*::::::::"),
	(0,     0,     0,     'W',     14,     0, ":::::::*::::::::"),
	(1,     0,     0,     'W',     15,     0, ":::::::*::::::::"),
	(0,     0,     1,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     2,     0, ":::::::::B::::::"),
	(0,     0,     1,     'W',     0,     0, "::*::::::B::::::"),
	(0,     1,     0,     'W',     12,     0, "W:*::::::B::::::"),
	(0,     1,     1,     'B',     11,     1, "::::::::::::::::"),
	(0,     1,     0,     ':',     2,     0, ":::::::::::B::::"),
	(0,     0,     1,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     9,     0, ":::::::::B::::::"),
	(0,     0,     1,     '*',     9,     0, ":::::::::B::::::"),
	(0,     0,     1,     ':',     1,     0, ":::::::::W::::::"),
	(0,     0,     1,     '*',     12,     0, ":::::::::W::::::"),
	(0,     0,     0,     'B',     2,     0, ":::::::::W::*:::"),
	(0,     0,     1,     'W',     12,     0, ":::::::::W::*:::"),
	(0,     0,     1,     '*',     10,     0, ":::::::::W::W:::"),
	(0,     0,     0,     'W',     3,     0, ":::::::::W*:W:::"),
	(0,     0,     0,     '*',     2,     0, ":::::::::W*:W:::"),
	(0,     0,     0,     '*',     0,     0, ":::::::::W*:W:::"),
	(0,     0,     0,     '*',     0,     0, ":::::::::W*:W:::"),
	(0,     0,     0,     'W',     11,     0, ":::::::::W*:W:::"),
	(1,     0,     0,     'B',     14,     0, ":::::::::W*:W:::"),
	(0,     0,     0,     'B',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     12,     0, "::::::*:::::::::"),
	(0,     0,     1,     'W',     11,     0, "::::::*:::::::::"),
	(0,     0,     1,     '*',     2,     0, "::::::*::::W::::"),
	(0,     0,     0,     '*',     15,     0, "::*:::*::::W::::"),
	(0,     0,     0,     ':',     0,     0, "::*:::*::::W::::"),
	(0,     0,     0,     ':',     0,     0, "::*:::*::::W::::"),
	(0,     0,     0,     'B',     10,     0, "::*:::*::::W::::"),
	(0,     0,     0,     'W',     11,     0, "::*:::*::::W::::"),
	(0,     0,     0,     ':',     5,     0, "::*:::*::::W::::"),
	(0,     0,     0,     'B',     12,     0, "::*:::*::::W::::"),
	(0,     0,     0,     ':',     10,     0, "::*:::*::::W::::"),
	(0,     0,     0,     ':',     9,     0, "::*:::*::::W::::"),
	(0,     0,     0,     'W',     3,     0, "::*:::*::::W::::"),
	(0,     0,     0,     '*',     9,     0, "::*:::*::::W::::"),
	(0,     0,     0,     ':',     5,     0, "::*:::*::::W::::"),
	(0,     1,     1,     '*',     15,     0, "::*:::*::::W::::"),
	(0,     0,     1,     'B',     15,     0, ":::::::::::::::*"),
	(0,     0,     1,     ':',     13,     0, ":::::::::::::::B"),
	(0,     0,     1,     '*',     5,     0, ":::::::::::::::B"),
	(0,     0,     0,     'W',     15,     0, ":::::*:::::::::B"),
	(0,     0,     0,     ':',     13,     0, ":::::*:::::::::B"),
	(0,     0,     0,     '*',     4,     0, ":::::*:::::::::B"),
	(0,     0,     0,     'B',     10,     0, ":::::*:::::::::B"),
	(0,     0,     1,     'W',     0,     0, ":::::*:::::::::B"),
	(0,     0,     1,     '*',     2,     0, "W::::*:::::::::B"),
	(0,     0,     1,     '*',     13,     0, "W:*::*:::::::::B"),
	(0,     0,     0,     'B',     9,     0, "W:*::*:::::::*:B"),
	(0,     0,     1,     ':',     12,     0, "W:*::*:::::::*:B"),
	(0,     1,     0,     ':',     10,     0, "W:*::*:::::::*:B"),
	(0,     0,     0,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     12,     0, "W:::::::::::::::"),
	(0,     0,     1,     'B',     13,     0, "W:::::::::::::::"),
	(0,     0,     0,     ':',     10,     0, "W::::::::::::B::"),
	(0,     0,     0,     '*',     15,     0, "W::::::::::::B::"),
	(0,     0,     0,     'B',     1,     0, "W::::::::::::B::"),
	(0,     0,     1,     'W',     10,     0, "W::::::::::::B::"),
	(0,     1,     1,     'W',     3,     0, "W:::::::::W::B::"),
	(0,     0,     0,     '*',     8,     0, ":::W::::::::::::"),
	(0,     0,     0,     '*',     3,     0, ":::W::::::::::::"),
	(0,     0,     0,     ':',     12,     0, ":::W::::::::::::"),
	(0,     0,     1,     'W',     13,     0, ":::W::::::::::::"),
	(0,     0,     0,     'B',     6,     0, ":::W:::::::::W::"),
	(0,     0,     1,     ':',     12,     0, ":::W:::::::::W::"),
	(0,     0,     1,     '*',     7,     0, ":::W:::::::::W::"),
	(0,     0,     0,     '*',     13,     0, ":::W:::*:::::W::"),
	(0,     1,     0,     'B',     11,     0, ":::W:::*:::::W::"),
	(0,     1,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     0,     0, "::::::::::::::B:"),
	(0,     0,     0,     'B',     0,     0, "::::::::::::::B:"),
	(0,     0,     0,     '*',     0,     0, "::::::::::::::B:"),
	(0,     0,     0,     'B',     10,     0, "::::::::::::::B:"),
	(0,     0,     1,     'W',     2,     0, "::::::::::::::B:"),
	(0,     0,     0,     'B',     13,     0, "::W:::::::::::B:"),
	(0,     0,     0,     '*',     2,     0, "::W:::::::::::B:"),
	(0,     0,     0,     '*',     1,     0, "::W:::::::::::B:"),
	(0,     0,     1,     'W',     1,     0, "::W:::::::::::B:"),
	(0,     0,     0,     'B',     4,     0, ":WW:::::::::::B:"),
	(0,     0,     1,     'W',     8,     0, ":WW:::::::::::B:"),
	(0,     0,     0,     'W',     9,     0, ":WW:::::W:::::B:"),
	(0,     1,     0,     'W',     8,     0, ":WW:::::W:::::B:"),
	(0,     0,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     9,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     4,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     14,     0, "::::B:::::::::::"),
	(0,     0,     0,     '*',     3,     0, "::::::::::::::B:"),
	(0,     0,     0,     'B',     13,     0, "::::::::::::::B:"),
	(0,     0,     1,     'W',     6,     0, "::::::::::::::B:"),
	(0,     0,     0,     ':',     12,     0, "::::::W:::::::B:"),
	(1,     0,     0,     ':',     8,     0, "::::::W:::::::B:"),
	(0,     0,     0,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     13,     0, "::*:::::::::::::"),
	(0,     0,     1,     'B',     9,     0, "::*:::::::::::::"),
	(0,     0,     1,     ':',     9,     0, "::*::::::B::::::"),
	(0,     0,     0,     ':',     5,     0, "::*::::::B::::::"),
	(1,     0,     1,     'W',     2,     0, "::*::::::B::::::"),
	(0,     0,     0,     ':',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     15,     0, ":::::::B::::::::"),
	(0,     0,     0,     'W',     15,     0, ":::::::B:::::::W"),
	(0,     0,     1,     ':',     15,     0, ":::::::B:::::::W"),
	(0,     0,     0,     'B',     9,     0, ":::::::B:::::::W"),
	(0,     0,     0,     ':',     12,     0, ":::::::B:::::::W"),
	(0,     1,     1,     'B',     12,     0, ":::::::B:::::::W"),
	(0,     0,     1,     'W',     11,     0, "::::::::::::B:::"),
	(0,     0,     1,     ':',     15,     0, ":::::::::::WB:::"),
	(0,     0,     0,     'W',     4,     0, ":::::::::::WB:::"),
	(0,     0,     1,     'W',     9,     0, ":::::::::::WB:::"),
	(0,     0,     0,     '*',     15,     0, ":::::::::W:WB:::"),
	(0,     0,     0,     '*',     7,     0, ":::::::::W:WB:::"),
	(0,     0,     0,     'B',     12,     0, ":::::::::W:WB:::"),
	(0,     0,     0,     'W',     13,     0, ":::::::::W:WB:::"),
	(0,     0,     1,     '*',     13,     0, ":::::::::W:WB:::"),
	(0,     0,     0,     'B',     12,     0, ":::::::::W:WB*::"),
	(0,     0,     1,     'W',     8,     0, ":::::::::W:WB*::"),
	(0,     0,     0,     'W',     9,     0, "::::::::WW:WB*::"),
	(0,     0,     0,     ':',     1,     0, "::::::::WW:WB*::"),
	(0,     0,     1,     '*',     9,     0, "::::::::WW:WB*::"),
	(0,     0,     1,     'B',     6,     0, "::::::::WB:WB*::"),
	(0,     0,     1,     ':',     9,     0, "::::::B:WB:WB*::"),
	(0,     0,     0,     'W',     8,     0, "::::::B:WB:WB*::"),
	(0,     0,     1,     '*',     13,     0, "::::::B:WB:WB*::"),
	(0,     0,     0,     ':',     2,     0, "::::::B:WB:WB:::"),
	(0,     0,     0,     '*',     11,     0, "::::::B:WB:WB:::"),
	(0,     0,     1,     '*',     1,     0, "::::::B:WB:WB:::"),
	(0,     0,     0,     'W',     5,     0, ":*::::B:WB:WB:::"),
	(0,     0,     1,     '*',     4,     0, ":*::::B:WB:WB:::"),
	(0,     0,     0,     '*',     15,     0, ":*::*:B:WB:WB:::"),
	(0,     0,     0,     '*',     11,     0, ":*::*:B:WB:WB:::"),
	(0,     1,     1,     ':',     4,     0, ":*::*:B:WB:WB:::"),
	(0,     0,     1,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     4,     0, "W:::::::::::::::"),
	(0,     1,     1,     ':',     12,     0, "W:::W:::::::::::"),
	(0,     0,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     3,     1, "::::::::::::::::"),
	(0,     1,     1,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     0,     0, "::::::*:::::::::"),
	(0,     0,     1,     'B',     14,     0, "B:::::*:::::::::"),
	(0,     0,     0,     'W',     15,     0, "B:::::*:::::::B:"),
	(0,     0,     1,     'B',     2,     0, "B:::::*:::::::B:"),
	(0,     0,     1,     'B',     4,     0, "B:B:::*:::::::B:"),
	(0,     0,     1,     'W',     12,     0, "B:B:B:*:::::::B:"),
	(0,     0,     1,     ':',     7,     0, "B:B:B:*:::::W:B:"),
	(0,     0,     0,     'W',     13,     0, "B:B:B:*:::::W:B:"),
	(0,     0,     0,     'B',     15,     0, "B:B:B:*:::::W:B:"),
	(0,     1,     1,     ':',     12,     0, "B:B:B:*:::::W:B:"),
	(0,     0,     0,     'B',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     10,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     13,     0, "::::::::::B:::::"),
	(0,     0,     0,     ':',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     12,     0, ":::::::::::::B::"),
	(0,     0,     0,     ':',     14,     0, ":::::::::::::B::"),
	(0,     0,     0,     'B',     1,     0, ":::::::::::::B::"),
	(0,     0,     1,     'B',     11,     0, ":::::::::::::B::"),
	(0,     0,     0,     ':',     0,     0, ":::::::::::B:B::"),
	(0,     0,     0,     'W',     9,     0, ":::::::::::B:B::"),
	(0,     1,     0,     ':',     13,     0, ":::::::::::B:B::"),
	(0,     0,     1,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     11,     0, "::::::::::W:::::"),
	(0,     0,     0,     'B',     10,     0, "::::::::::W*::::"),
	(0,     0,     1,     'B',     0,     0, "::::::::::W*::::"),
	(0,     0,     1,     '*',     12,     0, "B:::::::::W*::::"),
	(0,     0,     1,     '*',     2,     0, "B:::::::::W**:::"),
	(0,     0,     0,     '*',     7,     0, "B:*:::::::W**:::"),
	(0,     0,     1,     '*',     1,     0, "B:*:::::::W**:::"),
	(0,     0,     1,     ':',     11,     0, "B**:::::::W**:::"),
	(0,     0,     1,     ':',     12,     0, "B**:::::::W**:::"),
	(0,     0,     0,     '*',     2,     0, "B**:::::::W**:::"),
	(0,     0,     0,     'B',     12,     0, "B**:::::::W**:::"),
	(0,     0,     1,     'B',     0,     0, "B**:::::::W**:::"),
	(0,     1,     1,     '*',     14,     0, "B**:::::::W**:::"),
	(0,     0,     0,     ':',     10,     0, "::::::::::::::*:"),
	(0,     0,     1,     'W',     4,     0, "::::::::::::::*:"),
	(0,     0,     1,     '*',     6,     0, "::::W:::::::::*:"),
	(0,     0,     1,     '*',     5,     0, "::::W:*:::::::*:"),
	(0,     0,     1,     'B',     11,     0, "::::W**:::::::*:"),
	(0,     0,     0,     ':',     15,     0, "::::W**::::B::*:"),
	(0,     0,     0,     '*',     0,     0, "::::W**::::B::*:"),
	(0,     0,     0,     'W',     8,     0, "::::W**::::B::*:"),
	(0,     0,     1,     '*',     2,     0, "::::W**::::B::*:"),
	(0,     0,     1,     'W',     15,     0, "::*:W**::::B::*:"),
	(0,     0,     1,     '*',     13,     0, "::*:W**::::B::*W"),
	(0,     0,     0,     ':',     10,     0, "::*:W**::::B:**W"),
	(0,     0,     1,     ':',     12,     0, "::*:W**::::B:**W"),
	(0,     0,     1,     'W',     2,     0, "::*:W**::::B:**W"),
	(0,     0,     1,     'B',     6,     0, "::W:W**::::B:**W"),
	(0,     1,     0,     'W',     0,     0, "::W:W*B::::B:**W"),
	(0,     0,     0,     '*',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     12,     1, "::::::::::::::::"),
	(0,     1,     1,     '*',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     6,     0, "::::::::*:::::::"),
	(0,     0,     0,     'B',     7,     0, "::::::::*:::::::"),
	(0,     0,     1,     '*',     3,     0, "::::::::*:::::::"),
	(0,     1,     0,     ':',     4,     0, ":::*::::*:::::::"),
	(0,     0,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     1,     1,     'W',     12,     0, "::::::::::::W:::"),
	(1,     0,     0,     '*',     5,     0, "::::::::::::W:::"),
	(0,     1,     1,     'B',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     10,     0, "B:::::::::::::::"),
	(0,     1,     1,     '*',     2,     0, "B:::::::::::::::"),
	(0,     1,     1,     '*',     1,     0, "::*:::::::::::::"),
	(0,     0,     0,     'B',     2,     0, ":*::::::::::::::"),
	(0,     0,     1,     'B',     11,     0, ":*::::::::::::::"),
	(0,     0,     0,     'W',     6,     0, ":*:::::::::B::::"),
	(0,     0,     0,     'B',     5,     0, ":*:::::::::B::::"),
	(0,     0,     1,     ':',     2,     0, ":*:::::::::B::::"),
	(0,     0,     1,     ':',     2,     0, ":*:::::::::B::::"),
	(0,     0,     1,     'B',     15,     0, ":*:::::::::B::::"),
	(0,     0,     0,     'B',     6,     0, ":*:::::::::B:::B"),
	(0,     0,     0,     ':',     13,     0, ":*:::::::::B:::B"),
	(0,     0,     0,     'B',     1,     0, ":*:::::::::B:::B"),
	(0,     0,     1,     'W',     13,     0, ":*:::::::::B:::B"),
	(0,     0,     1,     ':',     9,     0, ":*:::::::::B:W:B"),
	(0,     0,     0,     'W',     6,     0, ":*:::::::::B:W:B"),
	(0,     0,     0,     ':',     13,     0, ":*:::::::::B:W:B"),
	(0,     0,     0,     ':',     14,     0, ":*:::::::::B:W:B"),
	(0,     0,     1,     'B',     13,     0, ":*:::::::::B:W:B"),
	(0,     0,     1,     '*',     4,     0, ":*:::::::::B:B:B"),
	(0,     0,     0,     '*',     13,     0, ":*::*::::::B:B:B"),
	(0,     0,     0,     '*',     9,     0, ":*::*::::::B:B:B"),
	(0,     0,     1,     'W',     11,     0, ":*::*::::::B:B:B"),
	(0,     0,     1,     ':',     10,     0, ":*::*::::::W:B:B"),
	(0,     0,     1,     'B',     13,     0, ":*::*::::::W:B:B"),
	(0,     1,     1,     '*',     12,     0, ":*::*::::::W:B:B"),
	(0,     0,     1,     'W',     14,     0, "::::::::::::*:::"),
	(0,     1,     1,     ':',     1,     0, "::::::::::::*:W:"),
	(0,     0,     0,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     10,     0, ":::::::::::::B::"),
	(0,     0,     0,     'W',     9,     0, "::::::::::B::B::"),
	(0,     0,     1,     'B',     13,     0, "::::::::::B::B::"),
	(0,     0,     1,     ':',     3,     0, "::::::::::B::B::"),
	(0,     0,     1,     '*',     3,     0, "::::::::::B::B::"),
	(0,     0,     1,     'W',     15,     0, ":::*::::::B::B::"),
	(0,     0,     0,     ':',     15,     0, ":::*::::::B::B:W"),
	(0,     0,     1,     'B',     11,     0, ":::*::::::B::B:W"),
	(0,     0,     1,     '*',     5,     0, ":::*::::::BB:B:W"),
	(0,     0,     0,     ':',     13,     0, ":::*:*::::BB:B:W"),
	(0,     0,     0,     '*',     8,     0, ":::*:*::::BB:B:W"),
	(0,     1,     0,     ':',     0,     0, ":::*:*::::BB:B:W"),
	(0,     0,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     5,     0, "::::::::::*:::::"),
	(0,     0,     1,     '*',     3,     0, "::::::::::*:::::"),
	(0,     1,     0,     'B',     0,     0, ":::*::::::*:::::"),
	(0,     0,     1,     ':',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     1,     0, "*:::::::::::::::"),
	(0,     0,     1,     'W',     9,     0, "*W::::::::::::::"),
	(0,     0,     1,     'B',     7,     0, "*W:::::::W::::::"),
	(0,     0,     1,     'W',     2,     0, "*W:::::B:W::::::"),
	(0,     0,     1,     ':',     12,     0, "*WW::::B:W::::::"),
	(0,     0,     1,     ':',     11,     0, "*WW::::B:W::::::"),
	(0,     0,     1,     '*',     6,     0, "*WW::::B:W::::::"),
	(0,     0,     1,     '*',     7,     0, "*WW:::*B:W::::::"),
	(0,     0,     0,     ':',     0,     0, "*WW:::*W:W::::::"),
	(0,     0,     0,     ':',     9,     0, "*WW:::*W:W::::::"),
	(0,     0,     1,     'B',     5,     0, "*WW:::*W:W::::::"),
	(0,     0,     0,     '*',     12,     0, "*WW::B*W:W::::::"),
	(0,     0,     1,     '*',     1,     0, "*WW::B*W:W::::::"),
	(0,     0,     1,     'B',     8,     0, "*BW::B*W:W::::::"),
	(0,     0,     1,     '*',     1,     0, "*BW::B*WBW::::::"),
	(0,     0,     1,     ':',     6,     0, "*WW::B*WBW::::::"),
	(0,     0,     0,     'B',     4,     0, "*WW::B*WBW::::::"),
	(0,     1,     0,     ':',     3,     0, "*WW::B*WBW::::::"),
	(0,     0,     0,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     0,     0, ":::::::::::::::W"),
	(0,     0,     0,     ':',     6,     0, ":::::::::::::::W"),
	(0,     0,     0,     'W',     15,     0, ":::::::::::::::W"),
	(0,     0,     0,     'B',     2,     0, ":::::::::::::::W"),
	(0,     1,     1,     'B',     11,     0, ":::::::::::::::W"),
	(0,     0,     1,     'W',     4,     0, ":::::::::::B::::"),
	(0,     0,     1,     ':',     7,     0, "::::W::::::B::::"),
	(0,     0,     0,     'W',     1,     0, "::::W::::::B::::"),
	(0,     0,     1,     'B',     6,     0, "::::W::::::B::::"),
	(0,     0,     0,     'B',     12,     0, "::::W:B::::B::::"),
	(0,     1,     1,     ':',     11,     0, "::::W:B::::B::::"),
	(0,     0,     0,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     14,     0, ":::::B::::::::::"),
	(0,     0,     0,     '*',     7,     0, ":::::B::::::::::"),
	(0,     0,     1,     '*',     2,     0, ":::::B::::::::::"),
	(0,     0,     1,     '*',     12,     0, "::*::B::::::::::"),
	(0,     0,     0,     ':',     10,     0, "::*::B::::::*:::"),
	(1,     0,     1,     '*',     6,     0, "::*::B::::::*:::"),
	(0,     0,     1,     ':',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     15,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     9,     0, "::::::::::::B:::"),
	(0,     0,     1,     'W',     0,     0, "::::::::::::B:::"),
	(0,     1,     0,     'W',     3,     0, "W:::::::::::B:::"),
	(0,     0,     0,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     8,     0, "::::::W:::::::::"),
	(0,     0,     0,     'B',     7,     0, "::::::W:::::::::"),
	(0,     0,     0,     'B',     11,     0, "::::::W:::::::::"),
	(0,     0,     1,     'B',     9,     0, "::::::W:::::::::"),
	(0,     0,     1,     'W',     6,     0, "::::::W::B::::::"),
	(0,     0,     0,     ':',     3,     0, "::::::W::B::::::"),
	(0,     1,     0,     ':',     14,     0, "::::::W::B::::::"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     6,     0, "::::::W:::::::::"),
	(0,     0,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     4,     0, ":::::W::::::::::"),
	(0,     0,     0,     'W',     5,     0, "::::WW::::::::::"),
	(0,     0,     0,     'B',     3,     0, "::::WW::::::::::"),
	(0,     0,     0,     'B',     15,     0, "::::WW::::::::::"),
	(0,     0,     0,     ':',     1,     0, "::::WW::::::::::"),
	(0,     0,     0,     ':',     0,     0, "::::WW::::::::::"),
	(0,     0,     1,     'W',     11,     0, "::::WW::::::::::"),
	(0,     0,     1,     'B',     2,     0, "::::WW:::::W::::"),
	(0,     0,     1,     'B',     13,     0, "::B:WW:::::W::::"),
	(0,     0,     1,     '*',     7,     0, "::B:WW:::::W:B::"),
	(0,     0,     0,     '*',     14,     0, "::B:WW:*:::W:B::"),
	(0,     0,     0,     '*',     11,     0, "::B:WW:*:::W:B::"),
	(0,     0,     1,     'B',     10,     0, "::B:WW:*:::W:B::"),
	(0,     0,     1,     '*',     4,     0, "::B:WW:*::BW:B::"),
	(0,     0,     0,     ':',     10,     0, "::B:BW:*::BW:B::"),
	(0,     1,     1,     ':',     2,     0, "::B:BW:*::BW:B::"),
	(0,     0,     0,     '*',     5,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     6,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     2,     0, "::::::B:::::::::"),
	(0,     0,     1,     ':',     12,     0, "::::::B:::::::::"),
	(0,     0,     1,     ':',     6,     0, "::::::B:::::::::"),
	(0,     0,     1,     ':',     3,     0, "::::::B:::::::::"),
	(0,     0,     0,     '*',     13,     0, "::::::B:::::::::"),
	(0,     0,     1,     ':',     6,     0, "::::::B:::::::::"),
	(0,     0,     0,     'W',     3,     0, "::::::B:::::::::"),
	(0,     0,     0,     'W',     12,     0, "::::::B:::::::::"),
	(0,     0,     0,     '*',     13,     0, "::::::B:::::::::"),
	(0,     0,     0,     'B',     8,     0, "::::::B:::::::::"),
	(0,     0,     1,     'W',     11,     0, "::::::B:::::::::"),
	(0,     0,     1,     ':',     15,     0, "::::::B::::W::::"),
	(0,     0,     1,     'W',     15,     0, "::::::B::::W::::"),
	(0,     0,     1,     'B',     8,     0, "::::::B::::W:::W"),
	(0,     0,     1,     '*',     14,     0, "::::::B:B::W:::W"),
	(0,     0,     1,     'B',     3,     0, "::::::B:B::W::*W"),
	(0,     0,     0,     'B',     4,     0, ":::B::B:B::W::*W"),
	(0,     0,     0,     ':',     15,     0, ":::B::B:B::W::*W"),
	(0,     0,     1,     'B',     6,     0, ":::B::B:B::W::*W"),
	(0,     0,     1,     'B',     11,     0, ":::B::B:B::W::*W"),
	(0,     0,     1,     'W',     5,     0, ":::B::B:B::B::*W"),
	(0,     0,     0,     'B',     11,     0, ":::B:WB:B::B::*W"),
	(0,     0,     1,     ':',     0,     0, ":::B:WB:B::B::*W"),
	(0,     0,     0,     'B',     8,     0, ":::B:WB:B::B::*W"),
	(0,     0,     1,     'B',     9,     0, ":::B:WB:B::B::*W"),
	(0,     0,     0,     ':',     0,     0, ":::B:WB:BB:B::*W"),
	(0,     0,     0,     'W',     14,     0, ":::B:WB:BB:B::*W"),
	(0,     0,     0,     'B',     15,     0, ":::B:WB:BB:B::*W"),
	(0,     0,     1,     ':',     11,     0, ":::B:WB:BB:B::*W"),
	(0,     0,     1,     'W',     5,     0, ":::B:WB:BB:B::*W"),
	(0,     0,     0,     'B',     15,     0, ":::B:WB:BB:B::*W"),
	(0,     0,     1,     ':',     10,     0, ":::B:WB:BB:B::*W"),
	(0,     0,     1,     '*',     12,     0, ":::B:WB:BB:B::*W"),
	(0,     0,     0,     '*',     4,     0, ":::B:WB:BB:B*:*W"),
	(0,     0,     0,     'B',     13,     0, ":::B:WB:BB:B*:*W"),
	(0,     1,     0,     ':',     3,     0, ":::B:WB:BB:B*:*W"),
	(0,     0,     1,     ':',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     8,     1, "::::::::::::::::"),
	(0,     1,     0,     '*',     11,     0, "::::::::W:::::::"),
	(0,     0,     1,     'W',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     13,     0, "::::::W:::::::::"),
	(0,     0,     0,     'B',     15,     0, "::::::W:::::::::"),
	(0,     0,     1,     'W',     11,     0, "::::::W:::::::::"),
	(0,     1,     1,     'W',     11,     0, "::::::W::::W::::"),
	(0,     0,     1,     ':',     13,     0, ":::::::::::W::::"),
	(0,     0,     1,     'B',     4,     0, ":::::::::::W::::"),
	(0,     0,     0,     ':',     6,     0, "::::B::::::W::::"),
	(0,     0,     0,     'W',     4,     0, "::::B::::::W::::"),
	(0,     1,     1,     '*',     8,     0, "::::B::::::W::::"),
	(0,     1,     0,     'W',     15,     0, "::::::::*:::::::"),
	(0,     0,     0,     'W',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     2,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     4,     1, "::::::::::::::::"),
	(0,     1,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     7,     0, "::::::::::*:::::"),
	(0,     0,     1,     'W',     11,     0, "::::::::::*:::::"),
	(0,     0,     0,     'W',     1,     0, "::::::::::*W::::"),
	(0,     0,     1,     'B',     15,     0, "::::::::::*W::::"),
	(0,     0,     0,     'W',     9,     0, "::::::::::*W:::B"),
	(0,     0,     0,     'B',     13,     0, "::::::::::*W:::B"),
	(0,     0,     0,     ':',     2,     0, "::::::::::*W:::B"),
	(0,     0,     1,     'W',     0,     0, "::::::::::*W:::B"),
	(0,     0,     0,     'B',     1,     0, "W:::::::::*W:::B"),
	(0,     0,     0,     'B',     8,     0, "W:::::::::*W:::B"),
	(0,     0,     0,     'W',     6,     0, "W:::::::::*W:::B"),
	(0,     0,     0,     ':',     3,     0, "W:::::::::*W:::B"),
	(0,     0,     0,     'B',     5,     0, "W:::::::::*W:::B"),
	(0,     0,     1,     'B',     2,     0, "W:::::::::*W:::B"),
	(0,     0,     0,     '*',     2,     0, "W:B:::::::*W:::B"),
	(0,     0,     0,     ':',     11,     0, "W:B:::::::*W:::B"),
	(0,     0,     1,     'W',     6,     0, "W:B:::::::*W:::B"),
	(0,     0,     0,     'B',     7,     0, "W:B:::W:::*W:::B"),
	(0,     0,     1,     'W',     12,     0, "W:B:::W:::*W:::B"),
	(1,     0,     0,     ':',     6,     0, "W:B:::W:::*WW::B"),
	(0,     1,     0,     'W',     0,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     1,     1, "::::::::::::::::"),
	(0,     1,     1,     'B',     0,     0, ":W::::::::::::::"),
	(0,     0,     0,     'B',     13,     0, "B:::::::::::::::"),
	(0,     0,     1,     'W',     4,     0, "B:::::::::::::::"),
	(0,     0,     0,     '*',     11,     0, "B:::W:::::::::::"),
	(0,     0,     0,     ':',     5,     0, "B:::W:::::::::::"),
	(0,     0,     1,     'B',     9,     0, "B:::W:::::::::::"),
	(0,     0,     1,     'W',     8,     0, "B:::W::::B::::::"),
	(0,     0,     1,     '*',     11,     0, "B:::W:::WB::::::"),
	(0,     0,     0,     '*',     11,     0, "B:::W:::WB:*::::"),
	(0,     1,     0,     'B',     7,     0, "B:::W:::WB:*::::"),
	(0,     0,     1,     ':',     8,     1, "::::::::::::::::"),
	(0,     1,     0,     'B',     9,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     6,     0, ":::::*::::::::::"),
	(0,     0,     0,     'W',     11,     0, ":::::*W:::::::::"),
	(0,     0,     0,     ':',     12,     0, ":::::*W:::::::::"),
	(0,     0,     1,     'B',     14,     0, ":::::*W:::::::::"),
	(0,     0,     1,     ':',     7,     0, ":::::*W:::::::B:"),
	(0,     0,     0,     'B',     13,     0, ":::::*W:::::::B:"),
	(0,     0,     0,     '*',     7,     0, ":::::*W:::::::B:"),
	(0,     0,     1,     'W',     4,     0, ":::::*W:::::::B:"),
	(0,     0,     0,     'B',     7,     0, "::::W*W:::::::B:"),
	(0,     0,     1,     '*',     6,     0, "::::W*W:::::::B:"),
	(0,     0,     0,     ':',     6,     0, "::::W*B:::::::B:"),
	(0,     0,     0,     '*',     12,     0, "::::W*B:::::::B:"),
	(0,     0,     1,     '*',     5,     0, "::::W*B:::::::B:"),
	(0,     0,     0,     'B',     0,     0, "::::W:B:::::::B:"),
	(0,     0,     1,     '*',     6,     0, "::::W:B:::::::B:"),
	(0,     0,     0,     'B',     6,     0, "::::W:W:::::::B:"),
	(0,     0,     1,     ':',     14,     0, "::::W:W:::::::B:"),
	(0,     0,     1,     '*',     6,     0, "::::W:W:::::::B:"),
	(0,     0,     1,     'W',     12,     0, "::::W:B:::::::B:"),
	(0,     0,     0,     'W',     13,     0, "::::W:B:::::W:B:"),
	(0,     0,     0,     ':',     11,     0, "::::W:B:::::W:B:"),
	(0,     0,     0,     'W',     9,     0, "::::W:B:::::W:B:"),
	(0,     0,     0,     'B',     8,     0, "::::W:B:::::W:B:"),
	(0,     0,     1,     'W',     9,     0, "::::W:B:::::W:B:"),
	(0,     0,     1,     '*',     2,     0, "::::W:B::W::W:B:"),
	(0,     0,     0,     ':',     14,     0, "::*:W:B::W::W:B:"),
	(0,     0,     0,     ':',     9,     0, "::*:W:B::W::W:B:"),
	(0,     0,     0,     ':',     14,     0, "::*:W:B::W::W:B:"),
	(0,     0,     0,     'W',     12,     0, "::*:W:B::W::W:B:"),
	(0,     0,     1,     'B',     6,     0, "::*:W:B::W::W:B:"),
	(0,     0,     0,     ':',     15,     0, "::*:W:B::W::W:B:"),
	(0,     0,     0,     '*',     4,     0, "::*:W:B::W::W:B:"),
	(0,     0,     0,     'W',     1,     0, "::*:W:B::W::W:B:"),
	(0,     0,     0,     'W',     11,     0, "::*:W:B::W::W:B:"),
	(0,     0,     0,     'B',     2,     0, "::*:W:B::W::W:B:"),
	(0,     0,     0,     ':',     12,     0, "::*:W:B::W::W:B:"),
	(0,     0,     0,     'W',     0,     0, "::*:W:B::W::W:B:"),
	(0,     1,     1,     'W',     15,     0, "::*:W:B::W::W:B:"),
	(0,     0,     1,     'W',     5,     0, ":::::::::::::::W"),
	(0,     0,     0,     '*',     1,     0, ":::::W:::::::::W"),
	(0,     0,     1,     'B',     8,     0, ":::::W:::::::::W"),
	(0,     0,     0,     '*',     13,     0, ":::::W::B::::::W"),
	(0,     0,     0,     'W',     4,     0, ":::::W::B::::::W"),
	(0,     0,     0,     'B',     6,     0, ":::::W::B::::::W"),
	(0,     1,     0,     'B',     15,     0, ":::::W::B::::::W"),
	(0,     0,     0,     ':',     11,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     4,     0, "::::::::::::::*:"),
	(0,     0,     1,     ':',     7,     0, "::::::::::::::*:"),
	(0,     0,     0,     ':',     8,     0, "::::::::::::::*:"),
	(0,     0,     0,     'W',     4,     0, "::::::::::::::*:"),
	(0,     0,     1,     '*',     4,     0, "::::::::::::::*:"),
	(0,     0,     1,     'B',     14,     0, "::::*:::::::::*:"),
	(0,     1,     1,     'W',     13,     0, "::::*:::::::::B:"),
	(0,     0,     0,     'B',     11,     0, ":::::::::::::W::"),
	(0,     0,     1,     'W',     1,     0, ":::::::::::::W::"),
	(0,     0,     1,     ':',     2,     0, ":W:::::::::::W::"),
	(1,     0,     1,     ':',     4,     0, ":W:::::::::::W::"),
	(0,     0,     0,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     7,     1, "::::::::::::::::"),
	(1,     0,     0,     ':',     15,     0, ":::::::*::::::::"),
	(0,     0,     1,     'W',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     13,     0, ":::::::::::W::::"),
	(0,     0,     1,     'W',     4,     0, ":::::::::::W::::"),
	(0,     0,     1,     'B',     14,     0, "::::W::::::W::::"),
	(0,     0,     1,     ':',     14,     0, "::::W::::::W::B:"),
	(0,     1,     1,     '*',     6,     0, "::::W::::::W::B:"),
	(0,     0,     0,     ':',     8,     0, "::::::*:::::::::"),
	(0,     0,     0,     'W',     11,     0, "::::::*:::::::::"),
	(0,     0,     0,     'W',     7,     0, "::::::*:::::::::"),
	(0,     0,     0,     ':',     8,     0, "::::::*:::::::::"),
	(0,     0,     1,     ':',     4,     0, "::::::*:::::::::"),
	(0,     0,     1,     '*',     4,     0, "::::::*:::::::::"),
	(0,     1,     1,     '*',     11,     0, "::::*:*:::::::::"),
	(0,     0,     0,     '*',     11,     0, ":::::::::::*::::"),
	(0,     0,     1,     ':',     15,     0, ":::::::::::*::::"),
	(0,     0,     1,     'B',     1,     0, ":::::::::::*::::"),
	(0,     0,     1,     'B',     10,     0, ":B:::::::::*::::"),
	(0,     0,     1,     'B',     13,     0, ":B::::::::B*::::"),
	(0,     1,     1,     ':',     8,     0, ":B::::::::B*:B::"),
	(0,     0,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     6,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     7,     0, "::::*:::::::::::"),
	(0,     0,     1,     '*',     4,     0, "::::*:::::::::::"),
	(0,     0,     1,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     8,     0, "::::::::::::::*:"),
	(0,     0,     1,     'W',     6,     0, "::::::::::::::*:"),
	(0,     0,     1,     '*',     11,     0, "::::::W:::::::*:"),
	(0,     0,     0,     '*',     7,     0, "::::::W::::*::*:"),
	(0,     0,     1,     'W',     7,     0, "::::::W::::*::*:"),
	(0,     0,     0,     ':',     6,     0, "::::::WW:::*::*:"),
	(0,     0,     0,     'B',     12,     0, "::::::WW:::*::*:"),
	(0,     0,     1,     '*',     7,     0, "::::::WW:::*::*:"),
	(0,     0,     0,     'B',     5,     0, "::::::WB:::*::*:"),
	(0,     0,     0,     ':',     15,     0, "::::::WB:::*::*:"),
	(0,     0,     0,     'B',     8,     0, "::::::WB:::*::*:"),
	(0,     0,     0,     'W',     8,     0, "::::::WB:::*::*:"),
	(0,     0,     0,     'W',     6,     0, "::::::WB:::*::*:"),
	(0,     0,     1,     ':',     14,     0, "::::::WB:::*::*:"),
	(0,     0,     0,     '*',     2,     0, "::::::WB:::*::*:"),
	(0,     0,     0,     ':',     15,     0, "::::::WB:::*::*:"),
	(0,     0,     0,     '*',     11,     0, "::::::WB:::*::*:"),
	(0,     1,     1,     'W',     6,     0, "::::::WB:::*::*:"),
	(0,     0,     1,     'W',     14,     0, "::::::W:::::::::"),
	(0,     0,     0,     ':',     6,     0, "::::::W:::::::W:"),
	(0,     1,     1,     '*',     15,     0, "::::::W:::::::W:"),
	(0,     1,     1,     '*',     5,     0, ":::::::::::::::*"),
	(0,     0,     1,     'W',     3,     0, ":::::*::::::::::"),
	(0,     0,     0,     '*',     13,     0, ":::W:*::::::::::"),
	(0,     1,     0,     'W',     4,     0, ":::W:*::::::::::"),
	(0,     0,     1,     ':',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     4,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     2,     0, ":::::W::::::::::"),
	(0,     0,     0,     'W',     9,     0, ":::::W::::::::::"),
	(0,     0,     0,     ':',     7,     0, ":::::W::::::::::"),
	(0,     0,     0,     '*',     10,     0, ":::::W::::::::::"),
	(0,     1,     1,     'W',     3,     0, ":::::W::::::::::"),
	(0,     0,     1,     ':',     3,     0, ":::W::::::::::::"),
	(0,     0,     1,     '*',     7,     0, ":::W::::::::::::"),
	(0,     0,     0,     'B',     12,     0, ":::W:::*::::::::"),
	(0,     0,     1,     'W',     15,     0, ":::W:::*::::::::"),
	(0,     0,     1,     'W',     4,     0, ":::W:::*:::::::W"),
	(0,     0,     1,     '*',     9,     0, ":::WW::*:::::::W"),
	(0,     0,     0,     ':',     7,     0, ":::WW::*:*:::::W"),
	(0,     0,     0,     ':',     5,     0, ":::WW::*:*:::::W"),
	(0,     0,     0,     ':',     7,     0, ":::WW::*:*:::::W"),
	(0,     1,     1,     'B',     12,     0, ":::WW::*:*:::::W"),
	(0,     0,     0,     '*',     10,     0, "::::::::::::B:::"),
	(0,     0,     1,     'W',     3,     0, "::::::::::::B:::"),
	(1,     0,     1,     ':',     6,     0, ":::W::::::::B:::"),
	(0,     0,     0,     'B',     12,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     4,     0, "::::::::::::W:::"),
	(0,     1,     0,     '*',     6,     0, "::::::::::::W:::"),
	(0,     0,     1,     '*',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     8,     0, "::::::::*:::::::"),
	(0,     0,     1,     '*',     11,     0, "::::::::*:::::::"),
	(0,     0,     1,     ':',     14,     0, "::::::::*::*::::"),
	(0,     0,     1,     'W',     7,     0, "::::::::*::*::::"),
	(0,     0,     0,     'W',     6,     0, ":::::::W*::*::::"),
	(0,     1,     0,     '*',     13,     0, ":::::::W*::*::::"),
	(0,     0,     1,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     15,     0, ":::::*::::::::::"),
	(0,     0,     1,     'W',     14,     0, ":::::*::::::::::"),
	(0,     1,     0,     '*',     3,     0, ":::::*::::::::W:"),
	(0,     0,     1,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     8,     0, ":::B::::::::::::"),
	(0,     0,     1,     'W',     14,     0, ":::B::::*:::::::"),
	(0,     0,     1,     '*',     4,     0, ":::B::::*:::::W:"),
	(0,     0,     1,     ':',     0,     0, ":::B*:::*:::::W:"),
	(0,     0,     0,     '*',     15,     0, ":::B*:::*:::::W:"),
	(0,     0,     1,     'B',     5,     0, ":::B*:::*:::::W:"),
	(0,     0,     0,     'W',     3,     0, ":::B*B::*:::::W:"),
	(0,     1,     1,     '*',     1,     0, ":::B*B::*:::::W:"),
	(0,     0,     0,     ':',     1,     0, ":*::::::::::::::"),
	(0,     0,     1,     ':',     2,     0, ":*::::::::::::::"),
	(0,     0,     0,     ':',     15,     0, ":*::::::::::::::"),
	(0,     0,     0,     'B',     14,     0, ":*::::::::::::::"),
	(0,     0,     0,     'B',     1,     0, ":*::::::::::::::"),
	(0,     0,     1,     ':',     4,     0, ":*::::::::::::::"),
	(0,     0,     0,     ':',     0,     0, ":*::::::::::::::"),
	(1,     0,     1,     'B',     2,     0, ":*::::::::::::::"),
	(0,     0,     1,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     14,     0, ":::::::W::::::::"),
	(0,     0,     0,     ':',     15,     0, ":::::::W::::::::"),
	(0,     0,     1,     'B',     10,     0, ":::::::W::::::::"),
	(0,     0,     1,     'W',     5,     0, ":::::::W::B:::::"),
	(0,     0,     0,     ':',     14,     0, ":::::W:W::B:::::"),
	(0,     0,     0,     '*',     13,     0, ":::::W:W::B:::::"),
	(0,     0,     1,     'W',     5,     0, ":::::W:W::B:::::"),
	(0,     0,     1,     'B',     3,     0, ":::::W:W::B:::::"),
	(0,     0,     1,     'W',     15,     0, ":::B:W:W::B:::::"),
	(0,     0,     0,     'B',     11,     0, ":::B:W:W::B::::W"),
	(0,     0,     1,     'W',     1,     0, ":::B:W:W::B::::W"),
	(0,     0,     0,     '*',     14,     0, ":W:B:W:W::B::::W"),
	(0,     0,     0,     'W',     4,     0, ":W:B:W:W::B::::W"),
	(0,     0,     1,     '*',     15,     0, ":W:B:W:W::B::::W"),
	(0,     0,     0,     ':',     5,     0, ":W:B:W:W::B::::B"),
	(0,     0,     0,     ':',     3,     0, ":W:B:W:W::B::::B"),
	(0,     0,     1,     '*',     13,     0, ":W:B:W:W::B::::B"),
	(0,     0,     0,     'B',     3,     0, ":W:B:W:W::B::*:B"),
	(0,     0,     1,     'W',     13,     0, ":W:B:W:W::B::*:B"),
	(0,     0,     0,     'W',     3,     0, ":W:B:W:W::B::W:B"),
	(0,     0,     1,     'B',     1,     0, ":W:B:W:W::B::W:B"),
	(0,     0,     0,     'W',     12,     0, ":B:B:W:W::B::W:B"),
	(0,     0,     1,     'W',     1,     0, ":B:B:W:W::B::W:B"),
	(0,     0,     1,     'B',     10,     0, ":W:B:W:W::B::W:B"),
	(0,     0,     0,     ':',     3,     0, ":W:B:W:W::B::W:B"),
	(0,     0,     0,     '*',     3,     0, ":W:B:W:W::B::W:B"),
	(0,     0,     1,     'B',     12,     0, ":W:B:W:W::B::W:B"),
	(0,     0,     1,     'B',     14,     0, ":W:B:W:W::B:BW:B"),
	(0,     0,     1,     'B',     14,     0, ":W:B:W:W::B:BWBB"),
	(0,     0,     1,     ':',     3,     0, ":W:B:W:W::B:BWBB"),
	(0,     0,     1,     '*',     4,     0, ":W:B:W:W::B:BWBB"),
	(0,     0,     1,     '*',     2,     0, ":W:B*W:W::B:BWBB"),
	(0,     0,     0,     '*',     3,     0, ":W*B*W:W::B:BWBB"),
	(0,     0,     0,     ':',     3,     0, ":W*B*W:W::B:BWBB"),
	(0,     0,     0,     ':',     13,     0, ":W*B*W:W::B:BWBB"),
	(0,     0,     0,     'W',     7,     0, ":W*B*W:W::B:BWBB"),
	(0,     0,     0,     ':',     12,     0, ":W*B*W:W::B:BWBB"),
	(0,     0,     0,     ':',     6,     0, ":W*B*W:W::B:BWBB"),
	(0,     0,     1,     ':',     9,     0, ":W*B*W:W::B:BWBB"),
	(0,     0,     1,     ':',     12,     0, ":W*B*W:W::B:BWBB"),
	(0,     0,     0,     '*',     14,     0, ":W*B*W:W::B:BWBB"),
	(0,     0,     0,     'B',     9,     0, ":W*B*W:W::B:BWBB"),
	(0,     1,     0,     '*',     15,     0, ":W*B*W:W::B:BWBB"),
	(0,     0,     1,     'B',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     10,     0, ":::::::B::::::::"),
	(0,     0,     0,     ':',     15,     0, ":::::::B::B:::::"),
	(0,     1,     0,     '*',     1,     0, ":::::::B::B:::::"),
	(0,     0,     1,     'B',     11,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     15,     0, ":::::::::::B::::"),
	(0,     0,     0,     'W',     10,     0, ":::::::::::B::::"),
	(0,     0,     1,     'W',     14,     0, ":::::::::::B::::"),
	(0,     0,     0,     '*',     11,     0, ":::::::::::B::W:"),
	(0,     0,     0,     '*',     10,     0, ":::::::::::B::W:"),
	(0,     0,     0,     ':',     15,     0, ":::::::::::B::W:"),
	(0,     0,     1,     ':',     0,     0, ":::::::::::B::W:"),
	(0,     0,     0,     'W',     7,     0, ":::::::::::B::W:"),
	(0,     0,     1,     'B',     10,     0, ":::::::::::B::W:"),
	(0,     0,     1,     ':',     10,     0, "::::::::::BB::W:"),
	(0,     0,     0,     ':',     14,     0, "::::::::::BB::W:"),
	(0,     0,     1,     ':',     4,     0, "::::::::::BB::W:"),
	(0,     0,     0,     '*',     8,     0, "::::::::::BB::W:"),
	(0,     0,     1,     'B',     11,     0, "::::::::::BB::W:"),
	(0,     0,     0,     'W',     5,     0, "::::::::::BB::W:"),
	(0,     0,     0,     ':',     1,     0, "::::::::::BB::W:"),
	(0,     0,     1,     '*',     12,     0, "::::::::::BB::W:"),
	(0,     0,     0,     ':',     7,     0, "::::::::::BB*:W:"),
	(0,     1,     1,     'W',     2,     0, "::::::::::BB*:W:"),
	(0,     0,     1,     'B',     14,     0, "::W:::::::::::::"),
	(0,     0,     1,     '*',     14,     0, "::W:::::::::::B:"),
	(0,     0,     1,     '*',     11,     0, "::W:::::::::::W:"),
	(0,     0,     1,     '*',     1,     0, "::W::::::::*::W:"),
	(0,     0,     0,     'W',     15,     0, ":*W::::::::*::W:"),
	(0,     0,     1,     'B',     11,     0, ":*W::::::::*::W:"),
	(0,     0,     1,     'W',     15,     0, ":*W::::::::B::W:"),
	(0,     0,     0,     '*',     13,     0, ":*W::::::::B::WW"),
	(0,     1,     0,     'B',     11,     0, ":*W::::::::B::WW"),
	(0,     0,     1,     ':',     4,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     8,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     12,     0, "::::::::W:::::::"),
	(0,     0,     0,     'W',     10,     0, "::::::::W:::::::"),
	(0,     0,     1,     '*',     12,     0, "::::::::W:::::::"),
	(0,     0,     1,     'W',     12,     0, "::::::::W:::*:::"),
	(0,     0,     1,     ':',     4,     0, "::::::::W:::W:::"),
	(0,     0,     1,     'W',     4,     0, "::::::::W:::W:::"),
	(0,     0,     0,     '*',     3,     0, "::::W:::W:::W:::"),
	(0,     0,     0,     ':',     2,     0, "::::W:::W:::W:::"),
	(0,     1,     0,     'W',     7,     0, "::::W:::W:::W:::"),
	(0,     0,     1,     '*',     5,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     8,     0, ":::::*::::::::::"),
	(0,     0,     1,     '*',     13,     0, ":::::*::::::::::"),
	(0,     0,     0,     'W',     6,     0, ":::::*:::::::*::"),
	(0,     0,     1,     'B',     8,     0, ":::::*:::::::*::"),
	(0,     0,     1,     'W',     9,     0, ":::::*::B::::*::"),
	(0,     0,     1,     'B',     3,     0, ":::::*::BW:::*::"),
	(0,     1,     1,     '*',     7,     0, ":::B:*::BW:::*::"),
	(0,     0,     0,     'B',     14,     0, ":::::::*::::::::"),
	(0,     0,     0,     '*',     4,     0, ":::::::*::::::::"),
	(0,     0,     0,     'B',     0,     0, ":::::::*::::::::"),
	(0,     1,     0,     'W',     14,     0, ":::::::*::::::::"),
	(0,     0,     0,     ':',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     11,     0, "::::::::::*:::::"),
	(0,     0,     1,     'W',     15,     0, "::::::::::*:::::"),
	(0,     0,     1,     '*',     13,     0, "::::::::::*::::W"),
	(0,     0,     0,     'B',     14,     0, "::::::::::*::*:W"),
	(0,     1,     1,     '*',     10,     0, "::::::::::*::*:W"),
	(0,     0,     0,     ':',     11,     0, "::::::::::*:::::"),
	(0,     0,     0,     'B',     14,     0, "::::::::::*:::::"),
	(0,     0,     1,     '*',     8,     0, "::::::::::*:::::"),
	(0,     0,     0,     ':',     14,     0, "::::::::*:*:::::"),
	(0,     0,     0,     'B',     12,     0, "::::::::*:*:::::"),
	(0,     0,     0,     ':',     0,     0, "::::::::*:*:::::"),
	(0,     0,     1,     ':',     11,     0, "::::::::*:*:::::"),
	(0,     0,     1,     'B',     15,     0, "::::::::*:*:::::"),
	(0,     0,     1,     ':',     1,     0, "::::::::*:*::::B"),
	(0,     0,     1,     'W',     3,     0, "::::::::*:*::::B"),
	(0,     0,     0,     'B',     13,     0, ":::W::::*:*::::B"),
	(0,     0,     0,     '*',     4,     0, ":::W::::*:*::::B"),
	(0,     0,     0,     'B',     7,     0, ":::W::::*:*::::B"),
	(0,     0,     0,     'B',     8,     0, ":::W::::*:*::::B"),
	(0,     0,     1,     '*',     8,     0, ":::W::::*:*::::B"),
	(0,     0,     1,     'W',     0,     0, ":::W::::::*::::B"),
	(0,     1,     0,     ':',     14,     0, "W::W::::::*::::B"),
	(0,     0,     0,     'W',     9,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     12,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     3,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     15,     0, ":::B::::::::::::"),
	(0,     0,     1,     'W',     15,     0, ":::B::::::::::::"),
	(0,     0,     1,     '*',     12,     0, ":::B:::::::::::W"),
	(0,     0,     0,     ':',     1,     0, ":::B::::::::*::W"),
	(0,     0,     0,     ':',     14,     0, ":::B::::::::*::W"),
	(0,     0,     0,     'W',     14,     0, ":::B::::::::*::W"),
	(0,     0,     1,     'B',     2,     0, ":::B::::::::*::W"),
	(0,     0,     1,     ':',     3,     0, "::BB::::::::*::W"),
	(0,     0,     1,     'W',     9,     0, "::BB::::::::*::W"),
	(0,     0,     0,     'B',     10,     0, "::BB:::::W::*::W"),
	(0,     0,     1,     ':',     0,     0, "::BB:::::W::*::W"),
	(0,     0,     1,     'W',     3,     0, "::BB:::::W::*::W"),
	(0,     0,     1,     'W',     7,     0, "::BW:::::W::*::W"),
	(0,     0,     0,     'W',     2,     0, "::BW:::W:W::*::W"),
	(0,     0,     1,     '*',     11,     0, "::BW:::W:W::*::W"),
	(0,     0,     1,     'W',     9,     0, "::BW:::W:W:**::W"),
	(0,     0,     1,     'B',     2,     0, "::BW:::W:W:**::W"),
	(0,     0,     1,     ':',     11,     0, "::BW:::W:W:**::W"),
	(0,     1,     1,     '*',     9,     0, "::BW:::W:W:**::W"),
	(0,     0,     0,     ':',     2,     0, ":::::::::*::::::"),
	(0,     0,     1,     'B',     13,     0, ":::::::::*::::::"),
	(0,     0,     1,     ':',     2,     0, ":::::::::*:::B::"),
	(0,     1,     0,     'W',     6,     0, ":::::::::*:::B::"),
	(0,     0,     0,     '*',     1,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     2,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     15,     0, "::W:::::::::::::"),
	(0,     0,     1,     'B',     5,     0, "::W::::::::::::W"),
	(0,     0,     1,     ':',     6,     0, "::W::B:::::::::W"),
	(0,     1,     0,     ':',     3,     0, "::W::B:::::::::W"),
	(0,     0,     1,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     11,     0, "::::::::::::::B:"),
	(0,     0,     0,     'B',     6,     0, ":::::::::::*::B:"),
	(0,     0,     0,     '*',     15,     0, ":::::::::::*::B:"),
	(0,     0,     0,     '*',     13,     0, ":::::::::::*::B:"),
	(0,     0,     1,     'B',     9,     0, ":::::::::::*::B:"),
	(0,     0,     1,     '*',     4,     0, ":::::::::B:*::B:"),
	(0,     0,     0,     'W',     8,     0, "::::*::::B:*::B:"),
	(0,     0,     0,     'B',     0,     0, "::::*::::B:*::B:"),
	(0,     0,     1,     ':',     10,     0, "::::*::::B:*::B:"),
	(0,     0,     1,     'W',     9,     0, "::::*::::B:*::B:"),
	(0,     0,     0,     'W',     0,     0, "::::*::::W:*::B:"),
	(0,     0,     1,     'B',     1,     0, "::::*::::W:*::B:"),
	(0,     0,     0,     'B',     14,     0, ":B::*::::W:*::B:"),
	(0,     0,     1,     '*',     11,     0, ":B::*::::W:*::B:"),
	(0,     0,     0,     '*',     9,     0, ":B::*::::W::::B:"),
	(0,     0,     1,     ':',     2,     0, ":B::*::::W::::B:"),
	(0,     0,     0,     'W',     1,     0, ":B::*::::W::::B:"),
	(0,     0,     1,     ':',     11,     0, ":B::*::::W::::B:"),
	(0,     0,     0,     'B',     15,     0, ":B::*::::W::::B:"),
	(0,     0,     1,     'B',     13,     0, ":B::*::::W::::B:"),
	(0,     0,     0,     'B',     7,     0, ":B::*::::W:::BB:"),
	(0,     0,     1,     'B',     9,     0, ":B::*::::W:::BB:"),
	(0,     0,     0,     'B',     13,     0, ":B::*::::B:::BB:"),
	(0,     1,     1,     ':',     2,     0, ":B::*::::B:::BB:"),
	(0,     0,     0,     'B',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     7,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     6,     0, ":::::::W::::::::"),
	(0,     0,     0,     '*',     8,     0, "::::::*W::::::::"),
	(0,     0,     1,     '*',     3,     0, "::::::*W::::::::"),
	(0,     0,     1,     ':',     14,     0, ":::*::*W::::::::"),
	(0,     0,     0,     '*',     14,     0, ":::*::*W::::::::"),
	(0,     0,     0,     'W',     13,     0, ":::*::*W::::::::"),
	(0,     0,     0,     'W',     13,     0, ":::*::*W::::::::"),
	(0,     0,     0,     ':',     2,     0, ":::*::*W::::::::"),
	(0,     0,     0,     'W',     2,     0, ":::*::*W::::::::"),
	(0,     0,     0,     '*',     0,     0, ":::*::*W::::::::"),
	(0,     0,     1,     '*',     11,     0, ":::*::*W::::::::"),
	(0,     0,     0,     '*',     3,     0, ":::*::*W:::*::::"),
	(0,     0,     1,     'B',     11,     0, ":::*::*W:::*::::"),
	(0,     0,     0,     'W',     11,     0, ":::*::*W:::B::::"),
	(0,     0,     0,     'B',     2,     0, ":::*::*W:::B::::"),
	(0,     0,     0,     '*',     0,     0, ":::*::*W:::B::::"),
	(0,     0,     1,     'W',     5,     0, ":::*::*W:::B::::"),
	(0,     0,     0,     'B',     9,     0, ":::*:W*W:::B::::"),
	(0,     0,     1,     '*',     0,     0, ":::*:W*W:::B::::"),
	(0,     0,     0,     '*',     13,     0, "*::*:W*W:::B::::"),
	(0,     0,     0,     'W',     10,     0, "*::*:W*W:::B::::"),
	(0,     0,     0,     '*',     4,     0, "*::*:W*W:::B::::"),
	(0,     0,     0,     ':',     1,     0, "*::*:W*W:::B::::"),
	(0,     0,     0,     'W',     8,     0, "*::*:W*W:::B::::"),
	(0,     0,     0,     'B',     1,     0, "*::*:W*W:::B::::"),
	(0,     0,     1,     'W',     3,     0, "*::*:W*W:::B::::"),
	(0,     0,     0,     '*',     3,     0, "*::W:W*W:::B::::"),
	(0,     0,     0,     'B',     0,     0, "*::W:W*W:::B::::"),
	(0,     0,     0,     ':',     12,     0, "*::W:W*W:::B::::"),
	(0,     0,     1,     '*',     2,     0, "*::W:W*W:::B::::"),
	(0,     0,     0,     'B',     0,     0, "*:*W:W*W:::B::::"),
	(0,     0,     1,     'W',     2,     0, "*:*W:W*W:::B::::"),
	(0,     0,     0,     'B',     7,     0, "*:WW:W*W:::B::::"),
	(0,     0,     0,     'W',     12,     0, "*:WW:W*W:::B::::"),
	(0,     0,     0,     ':',     7,     0, "*:WW:W*W:::B::::"),
	(0,     0,     1,     'W',     7,     0, "*:WW:W*W:::B::::"),
	(0,     0,     1,     '*',     7,     0, "*:WW:W*W:::B::::"),
	(0,     0,     1,     'W',     11,     0, "*:WW:W*B:::B::::"),
	(0,     0,     0,     'B',     2,     0, "*:WW:W*B:::W::::"),
	(0,     0,     0,     'B',     7,     0, "*:WW:W*B:::W::::"),
	(0,     0,     0,     '*',     15,     0, "*:WW:W*B:::W::::"),
	(0,     0,     1,     'B',     8,     0, "*:WW:W*B:::W::::"),
	(0,     0,     0,     '*',     2,     0, "*:WW:W*BB::W::::"),
	(0,     0,     1,     'W',     12,     0, "*:WW:W*BB::W::::"),
	(0,     0,     0,     'B',     4,     0, "*:WW:W*BB::WW:::"),
	(0,     0,     0,     'B',     5,     0, "*:WW:W*BB::WW:::"),
	(0,     0,     1,     ':',     9,     0, "*:WW:W*BB::WW:::"),
	(0,     0,     1,     ':',     3,     0, "*:WW:W*BB::WW:::"),
	(0,     0,     1,     'B',     5,     0, "*:WW:W*BB::WW:::"),
	(0,     1,     0,     '*',     5,     0, "*:WW:B*BB::WW:::"),
	(0,     0,     0,     ':',     8,     1, "::::::::::::::::"),
	(0,     0,     1,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     'W',     14,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     12,     0, "::::::::::::::W:"),
	(0,     0,     1,     'W',     5,     0, "::::::::::::*:W:"),
	(0,     1,     0,     '*',     4,     0, ":::::W::::::*:W:"),
	(0,     0,     1,     'B',     1,     1, "::::::::::::::::"),
	(0,     0,     0,     'B',     11,     0, ":B::::::::::::::"),
	(0,     0,     1,     ':',     4,     0, ":B::::::::::::::"),
	(0,     0,     1,     'B',     11,     0, ":B::::::::::::::"),
	(0,     0,     0,     'B',     0,     0, ":B:::::::::B::::"),
	(0,     0,     0,     'W',     0,     0, ":B:::::::::B::::"),
	(0,     0,     1,     ':',     6,     0, ":B:::::::::B::::"),
	(0,     0,     1,     ':',     3,     0, ":B:::::::::B::::"),
	(0,     0,     0,     ':',     15,     0, ":B:::::::::B::::"),
	(0,     0,     0,     'W',     1,     0, ":B:::::::::B::::"),
	(0,     0,     1,     'B',     1,     0, ":B:::::::::B::::"),
	(0,     0,     0,     'W',     12,     0, ":B:::::::::B::::"),
	(0,     0,     1,     'B',     12,     0, ":B:::::::::B::::"),
	(0,     0,     1,     'B',     14,     0, ":B:::::::::BB:::"),
	(0,     0,     1,     'B',     11,     0, ":B:::::::::BB:B:"),
	(0,     0,     1,     '*',     9,     0, ":B:::::::::BB:B:"),
	(0,     0,     0,     ':',     13,     0, ":B:::::::*:BB:B:"),
	(0,     0,     0,     'W',     10,     0, ":B:::::::*:BB:B:"),
	(0,     1,     0,     '*',     13,     0, ":B:::::::*:BB:B:"),
	(0,     0,     1,     '*',     14,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     0,     0, "::::::::::::::*:"),
	(0,     1,     0,     'B',     9,     0, "::::::::::::::*:"),
	(0,     0,     1,     '*',     0,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     11,     0, "*:::::::::::::::"),
	(0,     0,     1,     '*',     12,     0, "*:::::::::::::::"),
	(0,     0,     0,     '*',     13,     0, "*:::::::::::*:::"),
	(0,     0,     0,     'W',     2,     0, "*:::::::::::*:::"),
	(0,     0,     0,     'B',     6,     0, "*:::::::::::*:::"),
	(0,     0,     0,     ':',     8,     0, "*:::::::::::*:::"),
	(0,     0,     0,     '*',     6,     0, "*:::::::::::*:::"),
	(0,     0,     0,     'W',     15,     0, "*:::::::::::*:::"),
	(0,     0,     0,     '*',     0,     0, "*:::::::::::*:::"),
	(0,     0,     1,     'B',     15,     0, "*:::::::::::*:::"),
	(0,     0,     0,     ':',     14,     0, "*:::::::::::*::B"),
	(0,     0,     0,     ':',     12,     0, "*:::::::::::*::B"),
	(0,     0,     0,     '*',     6,     0, "*:::::::::::*::B"),
	(0,     0,     0,     '*',     12,     0, "*:::::::::::*::B"),
	(0,     0,     1,     'W',     1,     0, "*:::::::::::*::B"),
	(0,     0,     1,     ':',     5,     0, "*W::::::::::*::B"),
	(0,     0,     1,     ':',     15,     0, "*W::::::::::*::B"),
	(0,     0,     1,     'W',     8,     0, "*W::::::::::*::B"),
	(0,     0,     0,     ':',     1,     0, "*W::::::W:::*::B"),
	(0,     0,     1,     ':',     6,     0, "*W::::::W:::*::B"),
	(0,     0,     1,     'W',     7,     0, "*W::::::W:::*::B"),
	(0,     0,     1,     'B',     7,     0, "*W:::::WW:::*::B"),
	(0,     0,     1,     ':',     3,     0, "*W:::::BW:::*::B"),
	(0,     0,     0,     ':',     14,     0, "*W:::::BW:::*::B"),
	(0,     0,     1,     '*',     4,     0, "*W:::::BW:::*::B"),
	(0,     1,     0,     'B',     3,     0, "*W::*::BW:::*::B"),
	(0,     0,     1,     'W',     13,     1, "::::::::::::::::"),
	(0,     0,     0,     ':',     9,     0, ":::::::::::::W::"),
	(0,     0,     0,     '*',     7,     0, ":::::::::::::W::"),
	(0,     0,     0,     ':',     3,     0, ":::::::::::::W::"),
	(0,     0,     0,     'W',     12,     0, ":::::::::::::W::"),
	(0,     1,     1,     'W',     14,     0, ":::::::::::::W::"),
	(0,     0,     0,     'B',     13,     0, "::::::::::::::W:"),
	(0,     0,     1,     'B',     1,     0, "::::::::::::::W:"),
	(0,     1,     0,     '*',     2,     0, ":B::::::::::::W:"),
	(0,     0,     1,     ':',     5,     1, "::::::::::::::::"),
	(0,     0,     1,     '*',     10,     1, "::::::::::::::::"),
	(0,     0,     1,     'B',     15,     0, "::::::::::*:::::"),
	(0,     0,     0,     'B',     6,     0, "::::::::::*::::B"),
	(0,     0,     0,     'W',     13,     0, "::::::::::*::::B"),
	(0,     0,     0,     'B',     9,     0, "::::::::::*::::B"),
	(0,     1,     0,     'W',     0,     0, "::::::::::*::::B"),
	(0,     0,     1,     'W',     10,     1, "::::::::::::::::"),
	(0,     0,     0,     '*',     9,     0, "::::::::::W:::::"),
	(0,     0,     1,     '*',     3,     0, "::::::::::W:::::"),
	(0,     0,     0,     'B',     7,     0, ":::*::::::W:::::"),
	(0,     0,     1,     'W',     7,     0, ":::*::::::W:::::"),
	(0,     0,     1,     '*',     5,     0, ":::*:::W::W:::::"),
	(0,     0,     1,     ':',     15,     0, ":::*:*:W::W:::::"),
	(0,     0,     1,     'B',     0,     0, ":::*:*:W::W:::::"),
	(0,     0,     1,     'W',     15,     0, "B::*:*:W::W:::::"),
	(0,     0,     0,     'B',     2,     0, "B::*:*:W::W::::W"),
	(0,     0,     1,     ':',     15,     0, "B::*:*:W::W::::W"),
	(0,     1,     1,     'B',     4,     0, "B::*:*:W::W::::W"),
	(0,     0,     1,     'B',     15,     0, "::::B:::::::::::"),
	(0,     0,     1,     '*',     9,     0, "::::B::::::::::B"),
	(0,     0,     1,     ':',     5,     0, "::::B::::*:::::B"),
	(0,     1,     1,     '*',     14,     0, "::::B::::*:::::B"),
	(0,     0,     0,     'W',     5,     0, "::::::::::::::*:"),
	(0,     0,     0,     '*',     15,     0, "::::::::::::::*:"),
	(0,     0,     1,     'W',     9,     0, "::::::::::::::*:"),
	(0,     0,     1,     '*',     9,     0, ":::::::::W::::*:"),
	(0,     0,     1,     ':',     12,     0, ":::::::::B::::*:"),
	(0,     0,     0,     'B',     6,     0, ":::::::::B::::*:"),
	(0,     0,     1,     '*',     13,     0, ":::::::::B::::*:"),
	(0,     0,     1,     'W',     13,     0, ":::::::::B:::**:"),
	(0,     0,     1,     'B',     10,     0, ":::::::::B:::W*:"),
	(0,     0,     0,     '*',     14,     0, ":::::::::BB::W*:"),
	(0,     0,     0,     'B',     13,     0, ":::::::::BB::W*:"),
	(0,     0,     0,     ':',     3,     0, ":::::::::BB::W*:"),
	(0,     0,     1,     'W',     13,     0, ":::::::::BB::W*:"),
	(0,     0,     1,     'B',     10,     0, ":::::::::BB::W*:"),
	(0,     0,     1,     '*',     10,     0, ":::::::::BB::W*:"),
	(0,     0,     0,     ':',     10,     0, ":::::::::BW::W*:")
	);
END PACKAGE ex4_data_pak;
